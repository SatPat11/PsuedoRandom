magic
tech sky130A
magscale 1 2
timestamp 1750956218
<< nwell >>
rect 1066 2159 18898 17425
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 382 1844 19490 17672
<< metal2 >>
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
<< obsm2 >>
rect 386 856 19484 19145
rect 386 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 19484 856
<< metal3 >>
rect 0 19728 800 19848
rect 0 19048 800 19168
rect 0 18368 800 18488
rect 0 17688 800 17808
rect 0 17008 800 17128
rect 0 16328 800 16448
rect 0 15648 800 15768
rect 0 14968 800 15088
rect 0 14288 800 14408
rect 0 13608 800 13728
rect 0 12928 800 13048
rect 0 12248 800 12368
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 0 10208 800 10328
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
rect 0 7488 800 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 0 5448 800 5568
rect 0 4768 800 4888
rect 0 4088 800 4208
rect 0 3408 800 3528
rect 0 2728 800 2848
rect 0 2048 800 2168
rect 0 1368 800 1488
rect 0 688 800 808
rect 0 8 800 128
<< obsm3 >>
rect 880 19648 19399 19820
rect 381 19248 19399 19648
rect 880 18968 19399 19248
rect 381 18568 19399 18968
rect 880 18288 19399 18568
rect 381 17888 19399 18288
rect 880 17608 19399 17888
rect 381 17208 19399 17608
rect 880 16928 19399 17208
rect 381 16528 19399 16928
rect 880 16248 19399 16528
rect 381 15848 19399 16248
rect 880 15568 19399 15848
rect 381 15168 19399 15568
rect 880 14888 19399 15168
rect 381 14488 19399 14888
rect 880 14208 19399 14488
rect 381 13808 19399 14208
rect 880 13528 19399 13808
rect 381 13128 19399 13528
rect 880 12848 19399 13128
rect 381 12448 19399 12848
rect 880 12168 19399 12448
rect 381 11768 19399 12168
rect 880 11488 19399 11768
rect 381 11088 19399 11488
rect 880 10808 19399 11088
rect 381 10408 19399 10808
rect 880 10128 19399 10408
rect 381 9728 19399 10128
rect 880 9448 19399 9728
rect 381 9048 19399 9448
rect 880 8768 19399 9048
rect 381 8368 19399 8768
rect 880 8088 19399 8368
rect 381 7688 19399 8088
rect 880 7408 19399 7688
rect 381 7008 19399 7408
rect 880 6728 19399 7008
rect 381 6328 19399 6728
rect 880 6048 19399 6328
rect 381 5648 19399 6048
rect 880 5368 19399 5648
rect 381 4968 19399 5368
rect 880 4688 19399 4968
rect 381 4288 19399 4688
rect 880 4008 19399 4288
rect 381 3608 19399 4008
rect 880 3328 19399 3608
rect 381 2928 19399 3328
rect 880 2648 19399 2928
rect 381 2248 19399 2648
rect 880 1968 19399 2248
rect 381 1568 19399 1968
rect 880 1288 19399 1568
rect 381 888 19399 1288
rect 880 608 19399 888
rect 381 208 19399 608
rect 880 35 19399 208
<< metal4 >>
rect -1076 -4 -756 19588
rect -416 656 -96 18928
rect 3163 -4 3483 19588
rect 3823 -4 4143 19588
rect 7602 -4 7922 19588
rect 8262 -4 8582 19588
rect 12041 -4 12361 19588
rect 12701 -4 13021 19588
rect 16480 -4 16800 19588
rect 17140 -4 17460 19588
rect 20060 656 20380 18928
rect 20720 -4 21040 19588
<< obsm4 >>
rect 795 19668 17973 19821
rect 795 2891 3083 19668
rect 3563 2891 3743 19668
rect 4223 2891 7522 19668
rect 8002 2891 8182 19668
rect 8662 2891 11961 19668
rect 12441 2891 12621 19668
rect 13101 2891 16400 19668
rect 16880 2891 17060 19668
rect 17540 2891 17973 19668
<< metal5 >>
rect -1076 19268 21040 19588
rect -416 18608 20380 18928
rect -1076 16004 21040 16324
rect -1076 15344 21040 15664
rect -1076 12196 21040 12516
rect -1076 11536 21040 11856
rect -1076 8388 21040 8708
rect -1076 7728 21040 8048
rect -1076 4580 21040 4900
rect -1076 3920 21040 4240
rect -416 656 20380 976
rect -1076 -4 21040 316
<< labels >>
rlabel metal4 s -1076 -4 -756 19588 4 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -1076 -4 21040 316 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -1076 19268 21040 19588 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 20720 -4 21040 19588 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3823 -4 4143 19588 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8262 -4 8582 19588 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12701 -4 13021 19588 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17140 -4 17460 19588 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -1076 4580 21040 4900 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -1076 8388 21040 8708 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -1076 12196 21040 12516 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -1076 16004 21040 16324 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s -416 656 -96 18928 4 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -416 656 20380 976 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -416 18608 20380 18928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 20060 656 20380 18928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3163 -4 3483 19588 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7602 -4 7922 19588 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12041 -4 12361 19588 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16480 -4 16800 19588 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1076 3920 21040 4240 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1076 7728 21040 8048 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1076 11536 21040 11856 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1076 15344 21040 15664 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 19728 800 19848 6 clk
port 3 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 rst_n
port 4 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 s_axi_araddr[0]
port 5 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 s_axi_araddr[1]
port 6 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 s_axi_araddr[2]
port 7 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 s_axi_araddr[3]
port 8 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 s_axi_arready
port 9 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 s_axi_arvalid
port 10 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 s_axi_awaddr[0]
port 11 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 s_axi_awaddr[1]
port 12 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 s_axi_awaddr[2]
port 13 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 s_axi_awaddr[3]
port 14 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 s_axi_awready
port 15 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 s_axi_awvalid
port 16 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 s_axi_bready
port 17 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 s_axi_bresp[0]
port 18 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 s_axi_bresp[1]
port 19 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 s_axi_bvalid
port 20 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 s_axi_rdata[0]
port 21 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 s_axi_rdata[1]
port 22 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 s_axi_rdata[2]
port 23 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 s_axi_rdata[3]
port 24 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 s_axi_rdata[4]
port 25 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 s_axi_rdata[5]
port 26 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 s_axi_rdata[6]
port 27 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 s_axi_rdata[7]
port 28 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 s_axi_rready
port 29 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 s_axi_rvalid
port 30 nsew signal output
rlabel metal3 s 0 688 800 808 6 s_axi_wdata[0]
port 31 nsew signal input
rlabel metal3 s 0 8 800 128 6 s_axi_wdata[1]
port 32 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 s_axi_wdata[2]
port 33 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 s_axi_wdata[3]
port 34 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 s_axi_wdata[4]
port 35 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 s_axi_wdata[5]
port 36 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 s_axi_wdata[6]
port 37 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 s_axi_wdata[7]
port 38 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 s_axi_wready
port 39 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 s_axi_wvalid
port 40 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1692386
string GDS_FILE /openlane/designs/lfsr_axi_top/runs/RUN_2025.06.26_16.40.27/results/signoff/lfsr_axi_top.magic.gds
string GDS_START 430668
<< end >>

