module lfsr_axi_top (clk,
    rst_n,
    s_axi_arready,
    s_axi_arvalid,
    s_axi_awready,
    s_axi_awvalid,
    s_axi_bready,
    s_axi_bvalid,
    s_axi_rready,
    s_axi_rvalid,
    s_axi_wready,
    s_axi_wvalid,
    s_axi_araddr,
    s_axi_awaddr,
    s_axi_bresp,
    s_axi_rdata,
    s_axi_wdata);
 input clk;
 input rst_n;
 output s_axi_arready;
 input s_axi_arvalid;
 output s_axi_awready;
 input s_axi_awvalid;
 input s_axi_bready;
 output s_axi_bvalid;
 input s_axi_rready;
 output s_axi_rvalid;
 output s_axi_wready;
 input s_axi_wvalid;
 input [3:0] s_axi_araddr;
 input [3:0] s_axi_awaddr;
 output [1:0] s_axi_bresp;
 output [7:0] s_axi_rdata;
 input [7:0] s_axi_wdata;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire net42;
 wire \u_axi_slave.ctrl_reg[0] ;
 wire \u_axi_slave.ctrl_reg[1] ;
 wire \u_axi_slave.ctrl_reg[2] ;
 wire \u_axi_slave.ctrl_reg[3] ;
 wire \u_axi_slave.ctrl_reg[4] ;
 wire \u_axi_slave.ctrl_reg[5] ;
 wire \u_axi_slave.ctrl_reg[6] ;
 wire \u_axi_slave.ctrl_reg[7] ;
 wire \u_axi_slave.lfsr_data[0] ;
 wire \u_axi_slave.lfsr_data[1] ;
 wire \u_axi_slave.lfsr_data[2] ;
 wire \u_axi_slave.lfsr_data[3] ;
 wire \u_axi_slave.lfsr_data[4] ;
 wire \u_axi_slave.lfsr_data[5] ;
 wire \u_axi_slave.lfsr_data[6] ;
 wire \u_axi_slave.lfsr_data[7] ;
 wire \u_axi_slave.seed_reg[0] ;
 wire \u_axi_slave.seed_reg[1] ;
 wire \u_axi_slave.seed_reg[2] ;
 wire \u_axi_slave.seed_reg[3] ;
 wire \u_axi_slave.seed_reg[4] ;
 wire \u_axi_slave.seed_reg[5] ;
 wire \u_axi_slave.seed_reg[6] ;
 wire \u_axi_slave.seed_reg[7] ;
 wire \u_axi_slave.taps_reg[0] ;
 wire \u_axi_slave.taps_reg[1] ;
 wire \u_axi_slave.taps_reg[2] ;
 wire \u_axi_slave.taps_reg[3] ;
 wire \u_axi_slave.taps_reg[4] ;
 wire \u_axi_slave.taps_reg[5] ;
 wire \u_axi_slave.taps_reg[6] ;
 wire \u_axi_slave.taps_reg[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;

 sky130_fd_sc_hd__and3_2 _151_ (.A(net22),
    .B(net11),
    .C(net24),
    .X(_044_));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 _152_ (.A(_044_),
    .SLEEP(net10),
    .X(_045_));
 sky130_fd_sc_hd__nor2_2 _153_ (.A(net8),
    .B(net7),
    .Y(_046_));
 sky130_fd_sc_hd__and3_2 _154_ (.A(net9),
    .B(_045_),
    .C(_046_),
    .X(_047_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_4 _155_ (.A(_047_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _156_ (.A0(\u_axi_slave.seed_reg[0] ),
    .A1(net14),
    .S(_048_),
    .X(_049_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _157_ (.A(_049_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _158_ (.A0(\u_axi_slave.seed_reg[1] ),
    .A1(net15),
    .S(_048_),
    .X(_050_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _159_ (.A(_050_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _160_ (.A0(\u_axi_slave.seed_reg[2] ),
    .A1(net16),
    .S(_048_),
    .X(_051_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _161_ (.A(_051_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _162_ (.A0(\u_axi_slave.seed_reg[3] ),
    .A1(net17),
    .S(_048_),
    .X(_052_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _163_ (.A(_052_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _164_ (.A0(\u_axi_slave.seed_reg[4] ),
    .A1(net18),
    .S(_048_),
    .X(_053_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _165_ (.A(_053_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _166_ (.A0(\u_axi_slave.seed_reg[5] ),
    .A1(net19),
    .S(_048_),
    .X(_054_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _167_ (.A(_054_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _168_ (.A0(\u_axi_slave.seed_reg[6] ),
    .A1(net20),
    .S(_048_),
    .X(_055_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _169_ (.A(_055_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_2 _170_ (.A0(\u_axi_slave.seed_reg[7] ),
    .A1(net21),
    .S(_048_),
    .X(_056_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _171_ (.A(_056_),
    .X(_007_));
 sky130_fd_sc_hd__and3b_2 _172_ (.A_N(net9),
    .B(_045_),
    .C(_046_),
    .X(_057_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_4 _173_ (.A(_057_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _174_ (.A0(\u_axi_slave.ctrl_reg[0] ),
    .A1(net14),
    .S(_058_),
    .X(_059_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _175_ (.A(_059_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _176_ (.A0(\u_axi_slave.ctrl_reg[1] ),
    .A1(net15),
    .S(_058_),
    .X(_060_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _177_ (.A(_060_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _178_ (.A0(\u_axi_slave.ctrl_reg[2] ),
    .A1(net16),
    .S(_058_),
    .X(_061_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _179_ (.A(_061_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _180_ (.A0(\u_axi_slave.ctrl_reg[3] ),
    .A1(net17),
    .S(_058_),
    .X(_062_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _181_ (.A(_062_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _182_ (.A0(\u_axi_slave.ctrl_reg[4] ),
    .A1(net18),
    .S(_058_),
    .X(_063_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _183_ (.A(_063_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _184_ (.A0(\u_axi_slave.ctrl_reg[5] ),
    .A1(net19),
    .S(_058_),
    .X(_064_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _185_ (.A(_064_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _186_ (.A0(\u_axi_slave.ctrl_reg[6] ),
    .A1(net20),
    .S(_058_),
    .X(_065_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _187_ (.A(_065_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _188_ (.A0(\u_axi_slave.ctrl_reg[7] ),
    .A1(net21),
    .S(_058_),
    .X(_066_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _189_ (.A(_066_),
    .X(_015_));
 sky130_fd_sc_hd__or2_0 _190_ (.A(net25),
    .B(_044_),
    .X(_067_));
 sky130_fd_sc_hd__a21boi_2 _191_ (.A1(net12),
    .A2(net25),
    .B1_N(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__buf_1 _192_ (.A(_068_),
    .X(_016_));
 sky130_fd_sc_hd__a21boi_2 _193_ (.A1(net22),
    .A2(net11),
    .B1_N(net24),
    .Y(_069_));
 sky130_fd_sc_hd__a21o_2 _194_ (.A1(net12),
    .A2(net25),
    .B1(_069_),
    .X(_017_));
 sky130_fd_sc_hd__nor2_2 _195_ (.A(\u_axi_slave.ctrl_reg[1] ),
    .B(\u_axi_slave.ctrl_reg[0] ),
    .Y(_070_));
 sky130_fd_sc_hd__and4_2 _196_ (.A(\u_axi_slave.lfsr_data[1] ),
    .B(\u_axi_slave.lfsr_data[0] ),
    .C(\u_axi_slave.taps_reg[0] ),
    .D(\u_axi_slave.taps_reg[1] ),
    .X(_071_));
 sky130_fd_sc_hd__a22oi_4 _197_ (.A1(\u_axi_slave.lfsr_data[0] ),
    .A2(\u_axi_slave.taps_reg[0] ),
    .B1(\u_axi_slave.taps_reg[1] ),
    .B2(\u_axi_slave.lfsr_data[1] ),
    .Y(_072_));
 sky130_fd_sc_hd__a22o_2 _198_ (.A1(\u_axi_slave.lfsr_data[4] ),
    .A2(\u_axi_slave.taps_reg[4] ),
    .B1(\u_axi_slave.taps_reg[5] ),
    .B2(\u_axi_slave.lfsr_data[5] ),
    .X(_073_));
 sky130_fd_sc_hd__nand4_4 _199_ (.A(\u_axi_slave.lfsr_data[5] ),
    .B(\u_axi_slave.lfsr_data[4] ),
    .C(\u_axi_slave.taps_reg[4] ),
    .D(\u_axi_slave.taps_reg[5] ),
    .Y(_074_));
 sky130_fd_sc_hd__o211a_2 _200_ (.A1(_071_),
    .A2(_072_),
    .B1(_073_),
    .C1(_074_),
    .X(_075_));
 sky130_fd_sc_hd__a211oi_4 _201_ (.A1(_073_),
    .A2(_074_),
    .B1(_071_),
    .C1(_072_),
    .Y(_076_));
 sky130_fd_sc_hd__a22o_2 _202_ (.A1(\u_axi_slave.lfsr_data[2] ),
    .A2(\u_axi_slave.taps_reg[2] ),
    .B1(\u_axi_slave.taps_reg[3] ),
    .B2(\u_axi_slave.lfsr_data[3] ),
    .X(_077_));
 sky130_fd_sc_hd__nand4_4 _203_ (.A(\u_axi_slave.lfsr_data[3] ),
    .B(\u_axi_slave.lfsr_data[2] ),
    .C(\u_axi_slave.taps_reg[2] ),
    .D(\u_axi_slave.taps_reg[3] ),
    .Y(_078_));
 sky130_fd_sc_hd__a22oi_4 _204_ (.A1(\u_axi_slave.lfsr_data[6] ),
    .A2(\u_axi_slave.taps_reg[6] ),
    .B1(\u_axi_slave.taps_reg[7] ),
    .B2(\u_axi_slave.lfsr_data[7] ),
    .Y(_079_));
 sky130_fd_sc_hd__and4_2 _205_ (.A(\u_axi_slave.lfsr_data[7] ),
    .B(\u_axi_slave.lfsr_data[6] ),
    .C(\u_axi_slave.taps_reg[6] ),
    .D(\u_axi_slave.taps_reg[7] ),
    .X(_080_));
 sky130_fd_sc_hd__a211o_2 _206_ (.A1(_077_),
    .A2(_078_),
    .B1(_079_),
    .C1(_080_),
    .X(_081_));
 sky130_fd_sc_hd__o211ai_4 _207_ (.A1(_079_),
    .A2(_080_),
    .B1(_077_),
    .C1(_078_),
    .Y(_082_));
 sky130_fd_sc_hd__o211a_2 _208_ (.A1(_075_),
    .A2(_076_),
    .B1(_081_),
    .C1(_082_),
    .X(_083_));
 sky130_fd_sc_hd__or4_2 _209_ (.A(\u_axi_slave.lfsr_data[5] ),
    .B(\u_axi_slave.lfsr_data[4] ),
    .C(\u_axi_slave.lfsr_data[7] ),
    .D(\u_axi_slave.lfsr_data[6] ),
    .X(_084_));
 sky130_fd_sc_hd__or4_2 _210_ (.A(\u_axi_slave.lfsr_data[1] ),
    .B(\u_axi_slave.lfsr_data[0] ),
    .C(\u_axi_slave.lfsr_data[3] ),
    .D(\u_axi_slave.lfsr_data[2] ),
    .X(_085_));
 sky130_fd_sc_hd__lpflow_clkinvkapwr_1 _211_ (.A(\u_axi_slave.ctrl_reg[1] ),
    .Y(_086_));
 sky130_fd_sc_hd__o21ai_2 _212_ (.A1(_084_),
    .A2(_085_),
    .B1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a211o_2 _213_ (.A1(_081_),
    .A2(_082_),
    .B1(_075_),
    .C1(_076_),
    .X(_088_));
 sky130_fd_sc_hd__or3b_2 _214_ (.A(_083_),
    .B(_087_),
    .C_N(_088_),
    .X(_089_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_8 _215_ (.A(_086_),
    .X(_090_));
 sky130_fd_sc_hd__or2_0 _216_ (.A(\u_axi_slave.ctrl_reg[1] ),
    .B(\u_axi_slave.ctrl_reg[0] ),
    .X(_091_));
 sky130_fd_sc_hd__buf_4 _217_ (.A(_091_),
    .X(_092_));
 sky130_fd_sc_hd__o21a_2 _218_ (.A1(_090_),
    .A2(\u_axi_slave.seed_reg[0] ),
    .B1(_092_),
    .X(_093_));
 sky130_fd_sc_hd__a22o_2 _219_ (.A1(\u_axi_slave.lfsr_data[0] ),
    .A2(_070_),
    .B1(_089_),
    .B2(_093_),
    .X(_018_));
 sky130_fd_sc_hd__nand2_4 _220_ (.A(_090_),
    .B(\u_axi_slave.ctrl_reg[0] ),
    .Y(_094_));
 sky130_fd_sc_hd__or2_0 _221_ (.A(\u_axi_slave.lfsr_data[1] ),
    .B(_092_),
    .X(_095_));
 sky130_fd_sc_hd__o221a_2 _222_ (.A1(_090_),
    .A2(\u_axi_slave.seed_reg[1] ),
    .B1(_094_),
    .B2(\u_axi_slave.lfsr_data[0] ),
    .C1(_095_),
    .X(_019_));
 sky130_fd_sc_hd__or2_0 _223_ (.A(\u_axi_slave.lfsr_data[2] ),
    .B(_092_),
    .X(_096_));
 sky130_fd_sc_hd__o221a_2 _224_ (.A1(_090_),
    .A2(\u_axi_slave.seed_reg[2] ),
    .B1(_094_),
    .B2(\u_axi_slave.lfsr_data[1] ),
    .C1(_096_),
    .X(_020_));
 sky130_fd_sc_hd__or3_2 _225_ (.A(\u_axi_slave.lfsr_data[2] ),
    .B(_070_),
    .C(_087_),
    .X(_097_));
 sky130_fd_sc_hd__o221a_2 _226_ (.A1(_090_),
    .A2(\u_axi_slave.seed_reg[3] ),
    .B1(_092_),
    .B2(\u_axi_slave.lfsr_data[3] ),
    .C1(_097_),
    .X(_021_));
 sky130_fd_sc_hd__or3_2 _227_ (.A(\u_axi_slave.lfsr_data[3] ),
    .B(_070_),
    .C(_087_),
    .X(_098_));
 sky130_fd_sc_hd__o221a_2 _228_ (.A1(_090_),
    .A2(\u_axi_slave.seed_reg[4] ),
    .B1(_092_),
    .B2(\u_axi_slave.lfsr_data[4] ),
    .C1(_098_),
    .X(_022_));
 sky130_fd_sc_hd__or2_0 _229_ (.A(\u_axi_slave.lfsr_data[5] ),
    .B(_092_),
    .X(_099_));
 sky130_fd_sc_hd__o221a_2 _230_ (.A1(_090_),
    .A2(\u_axi_slave.seed_reg[5] ),
    .B1(_094_),
    .B2(\u_axi_slave.lfsr_data[4] ),
    .C1(_099_),
    .X(_023_));
 sky130_fd_sc_hd__or2_0 _231_ (.A(\u_axi_slave.lfsr_data[6] ),
    .B(_092_),
    .X(_100_));
 sky130_fd_sc_hd__o221a_2 _232_ (.A1(_090_),
    .A2(\u_axi_slave.seed_reg[6] ),
    .B1(_094_),
    .B2(\u_axi_slave.lfsr_data[5] ),
    .C1(_100_),
    .X(_024_));
 sky130_fd_sc_hd__or2_0 _233_ (.A(\u_axi_slave.lfsr_data[7] ),
    .B(_092_),
    .X(_101_));
 sky130_fd_sc_hd__o221a_2 _234_ (.A1(_090_),
    .A2(\u_axi_slave.seed_reg[7] ),
    .B1(_094_),
    .B2(\u_axi_slave.lfsr_data[6] ),
    .C1(_101_),
    .X(_025_));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 _235_ (.A(net23),
    .SLEEP_B(net6),
    .X(_102_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_4 _236_ (.A(_102_),
    .X(_103_));
 sky130_fd_sc_hd__nand2_2 _237_ (.A(net13),
    .B(net34),
    .Y(_104_));
 sky130_fd_sc_hd__o21ai_0 _238_ (.A1(net34),
    .A2(_103_),
    .B1(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(_105_),
    .Y(_026_));
 sky130_fd_sc_hd__or3_4 _240_ (.A(net3),
    .B(net2),
    .C(net4),
    .X(_106_));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 _241_ (.A(net5),
    .SLEEP(_106_),
    .X(_107_));
 sky130_fd_sc_hd__or3b_4 _242_ (.A(net3),
    .B(net2),
    .C_N(net4),
    .X(_108_));
 sky130_fd_sc_hd__nor2_4 _243_ (.A(net5),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 _244_ (.A(\u_axi_slave.seed_reg[0] ),
    .SLEEP_B(_109_),
    .X(_110_));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 _245_ (.A(net5),
    .SLEEP(_108_),
    .X(_111_));
 sky130_fd_sc_hd__nor2_4 _246_ (.A(net5),
    .B(_106_),
    .Y(_112_));
 sky130_fd_sc_hd__a22o_2 _247_ (.A1(\u_axi_slave.lfsr_data[0] ),
    .A2(_111_),
    .B1(_112_),
    .B2(\u_axi_slave.ctrl_reg[0] ),
    .X(_113_));
 sky130_fd_sc_hd__nand2_4 _248_ (.A(net23),
    .B(net6),
    .Y(_114_));
 sky130_fd_sc_hd__a2111oi_2 _249_ (.A1(\u_axi_slave.taps_reg[0] ),
    .A2(_107_),
    .B1(_110_),
    .C1(_113_),
    .D1(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__o21ba_2 _250_ (.A1(net26),
    .A2(_103_),
    .B1_N(_115_),
    .X(_027_));
 sky130_fd_sc_hd__or4b_4 _251_ (.A(net3),
    .B(net2),
    .C(net4),
    .D_N(net5),
    .X(_116_));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 _252_ (.A(\u_axi_slave.taps_reg[1] ),
    .SLEEP(_116_),
    .X(_117_));
 sky130_fd_sc_hd__or2_0 _253_ (.A(net5),
    .B(_106_),
    .X(_118_));
 sky130_fd_sc_hd__o21ai_0 _254_ (.A1(_090_),
    .A2(_118_),
    .B1(_102_),
    .Y(_119_));
 sky130_fd_sc_hd__a22o_2 _255_ (.A1(\u_axi_slave.lfsr_data[1] ),
    .A2(_111_),
    .B1(_109_),
    .B2(\u_axi_slave.seed_reg[1] ),
    .X(_120_));
 sky130_fd_sc_hd__o32a_2 _256_ (.A1(_117_),
    .A2(_119_),
    .A3(_120_),
    .B1(_103_),
    .B2(net27),
    .X(_028_));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 _257_ (.A(\u_axi_slave.ctrl_reg[2] ),
    .SLEEP_B(_112_),
    .X(_121_));
 sky130_fd_sc_hd__lpflow_clkinvkapwr_1 _258_ (.A(\u_axi_slave.taps_reg[2] ),
    .Y(_122_));
 sky130_fd_sc_hd__o21ai_2 _259_ (.A1(_122_),
    .A2(_116_),
    .B1(_102_),
    .Y(_123_));
 sky130_fd_sc_hd__a221o_2 _260_ (.A1(\u_axi_slave.lfsr_data[2] ),
    .A2(_111_),
    .B1(_109_),
    .B2(\u_axi_slave.seed_reg[2] ),
    .C1(_123_),
    .X(_124_));
 sky130_fd_sc_hd__o22a_2 _261_ (.A1(net28),
    .A2(_103_),
    .B1(_121_),
    .B2(_124_),
    .X(_029_));
 sky130_fd_sc_hd__a22o_2 _262_ (.A1(\u_axi_slave.taps_reg[3] ),
    .A2(_107_),
    .B1(_109_),
    .B2(\u_axi_slave.seed_reg[3] ),
    .X(_125_));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 _263_ (.A(\u_axi_slave.lfsr_data[3] ),
    .SLEEP_B(_111_),
    .X(_126_));
 sky130_fd_sc_hd__a2111oi_2 _264_ (.A1(\u_axi_slave.ctrl_reg[3] ),
    .A2(_112_),
    .B1(_125_),
    .C1(_126_),
    .D1(_114_),
    .Y(_127_));
 sky130_fd_sc_hd__o21ba_2 _265_ (.A1(net29),
    .A2(_103_),
    .B1_N(_127_),
    .X(_030_));
 sky130_fd_sc_hd__lpflow_clkinvkapwr_1 _266_ (.A(\u_axi_slave.ctrl_reg[4] ),
    .Y(_128_));
 sky130_fd_sc_hd__o21ai_0 _267_ (.A1(_128_),
    .A2(_118_),
    .B1(_103_),
    .Y(_129_));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 _268_ (.A(\u_axi_slave.taps_reg[4] ),
    .SLEEP(_116_),
    .X(_130_));
 sky130_fd_sc_hd__a221o_2 _269_ (.A1(\u_axi_slave.lfsr_data[4] ),
    .A2(_111_),
    .B1(_109_),
    .B2(\u_axi_slave.seed_reg[4] ),
    .C1(_130_),
    .X(_131_));
 sky130_fd_sc_hd__o22a_2 _270_ (.A1(net30),
    .A2(_103_),
    .B1(_129_),
    .B2(_131_),
    .X(_031_));
 sky130_fd_sc_hd__a22o_2 _271_ (.A1(\u_axi_slave.taps_reg[5] ),
    .A2(_107_),
    .B1(_111_),
    .B2(\u_axi_slave.lfsr_data[5] ),
    .X(_132_));
 sky130_fd_sc_hd__a221o_2 _272_ (.A1(\u_axi_slave.seed_reg[5] ),
    .A2(_109_),
    .B1(_112_),
    .B2(\u_axi_slave.ctrl_reg[5] ),
    .C1(_114_),
    .X(_133_));
 sky130_fd_sc_hd__o22a_2 _273_ (.A1(net31),
    .A2(_103_),
    .B1(_132_),
    .B2(_133_),
    .X(_032_));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 _274_ (.A(\u_axi_slave.seed_reg[6] ),
    .SLEEP_B(_109_),
    .X(_134_));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 _275_ (.A(\u_axi_slave.lfsr_data[6] ),
    .SLEEP_B(_111_),
    .X(_135_));
 sky130_fd_sc_hd__a221o_2 _276_ (.A1(\u_axi_slave.taps_reg[6] ),
    .A2(_107_),
    .B1(_112_),
    .B2(\u_axi_slave.ctrl_reg[6] ),
    .C1(_114_),
    .X(_136_));
 sky130_fd_sc_hd__o32a_2 _277_ (.A1(_134_),
    .A2(_135_),
    .A3(_136_),
    .B1(_103_),
    .B2(net32),
    .X(_033_));
 sky130_fd_sc_hd__a22o_2 _278_ (.A1(\u_axi_slave.lfsr_data[7] ),
    .A2(_111_),
    .B1(_109_),
    .B2(\u_axi_slave.seed_reg[7] ),
    .X(_137_));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 _279_ (.A(\u_axi_slave.taps_reg[7] ),
    .SLEEP(_116_),
    .X(_138_));
 sky130_fd_sc_hd__a2111oi_2 _280_ (.A1(\u_axi_slave.ctrl_reg[7] ),
    .A2(_112_),
    .B1(_137_),
    .C1(_138_),
    .D1(_114_),
    .Y(_139_));
 sky130_fd_sc_hd__o21ba_2 _281_ (.A1(net33),
    .A2(_103_),
    .B1_N(_139_),
    .X(_034_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(net23),
    .Y(_140_));
 sky130_fd_sc_hd__o21ai_2 _283_ (.A1(_140_),
    .A2(net6),
    .B1(_104_),
    .Y(_035_));
 sky130_fd_sc_hd__and4b_2 _284_ (.A_N(net9),
    .B(net10),
    .C(_044_),
    .D(_046_),
    .X(_141_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_4 _285_ (.A(_141_),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _286_ (.A0(\u_axi_slave.taps_reg[0] ),
    .A1(net14),
    .S(_142_),
    .X(_143_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _287_ (.A(_143_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _288_ (.A0(\u_axi_slave.taps_reg[1] ),
    .A1(net15),
    .S(_142_),
    .X(_144_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _289_ (.A(_144_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _290_ (.A0(\u_axi_slave.taps_reg[2] ),
    .A1(net16),
    .S(_142_),
    .X(_145_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _291_ (.A(_145_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _292_ (.A0(\u_axi_slave.taps_reg[3] ),
    .A1(net17),
    .S(_142_),
    .X(_146_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _293_ (.A(_146_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(\u_axi_slave.taps_reg[4] ),
    .A1(net18),
    .S(_142_),
    .X(_147_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _295_ (.A(_147_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(\u_axi_slave.taps_reg[5] ),
    .A1(net19),
    .S(_142_),
    .X(_148_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _297_ (.A(_148_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _298_ (.A0(\u_axi_slave.taps_reg[6] ),
    .A1(net20),
    .S(_142_),
    .X(_149_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _299_ (.A(_149_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _300_ (.A0(\u_axi_slave.taps_reg[7] ),
    .A1(net21),
    .S(_142_),
    .X(_150_));
 sky130_fd_sc_hd__lpflow_clkbufkapwr_1 _301_ (.A(_150_),
    .X(_043_));
 sky130_fd_sc_hd__dfstp_2 _302_ (.CLK(clk),
    .D(_000_),
    .SET_B(net40),
    .Q(\u_axi_slave.seed_reg[0] ));
 sky130_fd_sc_hd__dfrtp_4 _303_ (.CLK(clk),
    .D(_001_),
    .RESET_B(net39),
    .Q(\u_axi_slave.seed_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _304_ (.CLK(clk),
    .D(_002_),
    .RESET_B(net36),
    .Q(\u_axi_slave.seed_reg[2] ));
 sky130_fd_sc_hd__dfstp_2 _305_ (.CLK(clk),
    .D(_003_),
    .SET_B(net39),
    .Q(\u_axi_slave.seed_reg[3] ));
 sky130_fd_sc_hd__dfstp_2 _306_ (.CLK(clk),
    .D(_004_),
    .SET_B(net37),
    .Q(\u_axi_slave.seed_reg[4] ));
 sky130_fd_sc_hd__dfrtp_4 _307_ (.CLK(clk),
    .D(_005_),
    .RESET_B(net39),
    .Q(\u_axi_slave.seed_reg[5] ));
 sky130_fd_sc_hd__dfrtp_4 _308_ (.CLK(clk),
    .D(_006_),
    .RESET_B(net37),
    .Q(\u_axi_slave.seed_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _309_ (.CLK(clk),
    .D(_007_),
    .RESET_B(net37),
    .Q(\u_axi_slave.seed_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _310_ (.CLK(clk),
    .D(_008_),
    .RESET_B(net39),
    .Q(\u_axi_slave.ctrl_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _311_ (.CLK(clk),
    .D(_009_),
    .RESET_B(net37),
    .Q(\u_axi_slave.ctrl_reg[1] ));
 sky130_fd_sc_hd__dfrtp_4 _312_ (.CLK(clk),
    .D(_010_),
    .RESET_B(net39),
    .Q(\u_axi_slave.ctrl_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _313_ (.CLK(clk),
    .D(_011_),
    .RESET_B(net37),
    .Q(\u_axi_slave.ctrl_reg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _314_ (.CLK(clk),
    .D(_012_),
    .RESET_B(net40),
    .Q(\u_axi_slave.ctrl_reg[4] ));
 sky130_fd_sc_hd__dfrtp_4 _315_ (.CLK(clk),
    .D(_013_),
    .RESET_B(net36),
    .Q(\u_axi_slave.ctrl_reg[5] ));
 sky130_fd_sc_hd__dfrtp_4 _316_ (.CLK(clk),
    .D(_014_),
    .RESET_B(net40),
    .Q(\u_axi_slave.ctrl_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _317_ (.CLK(clk),
    .D(_015_),
    .RESET_B(net39),
    .Q(\u_axi_slave.ctrl_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _318_ (.CLK(clk),
    .D(_016_),
    .RESET_B(net36),
    .Q(net25));
 sky130_fd_sc_hd__dfstp_2 _319_ (.CLK(clk),
    .D(_017_),
    .SET_B(net36),
    .Q(net24));
 sky130_fd_sc_hd__dfstp_4 _320_ (.CLK(clk),
    .D(_018_),
    .SET_B(net40),
    .Q(\u_axi_slave.lfsr_data[0] ));
 sky130_fd_sc_hd__dfrtp_2 _321_ (.CLK(clk),
    .D(_019_),
    .RESET_B(net36),
    .Q(\u_axi_slave.lfsr_data[1] ));
 sky130_fd_sc_hd__dfrtp_2 _322_ (.CLK(clk),
    .D(_020_),
    .RESET_B(net39),
    .Q(\u_axi_slave.lfsr_data[2] ));
 sky130_fd_sc_hd__dfstp_4 _323_ (.CLK(clk),
    .D(_021_),
    .SET_B(net37),
    .Q(\u_axi_slave.lfsr_data[3] ));
 sky130_fd_sc_hd__dfstp_4 _324_ (.CLK(clk),
    .D(_022_),
    .SET_B(net40),
    .Q(\u_axi_slave.lfsr_data[4] ));
 sky130_fd_sc_hd__dfrtp_2 _325_ (.CLK(clk),
    .D(_023_),
    .RESET_B(net39),
    .Q(\u_axi_slave.lfsr_data[5] ));
 sky130_fd_sc_hd__dfrtp_2 _326_ (.CLK(clk),
    .D(_024_),
    .RESET_B(net36),
    .Q(\u_axi_slave.lfsr_data[6] ));
 sky130_fd_sc_hd__dfrtp_2 _327_ (.CLK(clk),
    .D(_025_),
    .RESET_B(net40),
    .Q(\u_axi_slave.lfsr_data[7] ));
 sky130_fd_sc_hd__dfrtp_2 _328_ (.CLK(clk),
    .D(_026_),
    .RESET_B(net37),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_4 _329_ (.CLK(clk),
    .D(_027_),
    .RESET_B(net36),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_2 _330_ (.CLK(clk),
    .D(_028_),
    .RESET_B(net39),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_4 _331_ (.CLK(clk),
    .D(_029_),
    .RESET_B(net36),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_2 _332_ (.CLK(clk),
    .D(_030_),
    .RESET_B(net36),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_2 _333_ (.CLK(clk),
    .D(_031_),
    .RESET_B(net36),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_2 _334_ (.CLK(clk),
    .D(_032_),
    .RESET_B(net40),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_2 _335_ (.CLK(clk),
    .D(_033_),
    .RESET_B(net37),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_2 _336_ (.CLK(clk),
    .D(_034_),
    .RESET_B(net38),
    .Q(net33));
 sky130_fd_sc_hd__dfstp_4 _337_ (.CLK(clk),
    .D(_035_),
    .SET_B(net40),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_2 _338_ (.CLK(clk),
    .D(_036_),
    .RESET_B(net37),
    .Q(\u_axi_slave.taps_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _339_ (.CLK(clk),
    .D(_037_),
    .RESET_B(net1),
    .Q(\u_axi_slave.taps_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _340_ (.CLK(clk),
    .D(_038_),
    .RESET_B(net1),
    .Q(\u_axi_slave.taps_reg[2] ));
 sky130_fd_sc_hd__dfstp_2 _341_ (.CLK(clk),
    .D(_039_),
    .SET_B(net40),
    .Q(\u_axi_slave.taps_reg[3] ));
 sky130_fd_sc_hd__dfstp_2 _342_ (.CLK(clk),
    .D(_040_),
    .SET_B(net38),
    .Q(\u_axi_slave.taps_reg[4] ));
 sky130_fd_sc_hd__dfstp_2 _343_ (.CLK(clk),
    .D(_041_),
    .SET_B(net39),
    .Q(\u_axi_slave.taps_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _344_ (.CLK(clk),
    .D(_042_),
    .RESET_B(net38),
    .Q(\u_axi_slave.taps_reg[6] ));
 sky130_fd_sc_hd__dfstp_2 _345_ (.CLK(clk),
    .D(_043_),
    .SET_B(net37),
    .Q(\u_axi_slave.taps_reg[7] ));
 sky130_fd_sc_hd__conb_1 lfsr_axi_top_42 (.LO(net42));
 sky130_fd_sc_hd__buf_1 _348_ (.A(net24),
    .X(net35));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_145 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(s_axi_araddr[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(s_axi_araddr[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(s_axi_araddr[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(s_axi_araddr[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(s_axi_arvalid),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(s_axi_awaddr[0]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(s_axi_awaddr[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(s_axi_awaddr[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(s_axi_awaddr[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(s_axi_awvalid),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(s_axi_bready),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(s_axi_rready),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(s_axi_wdata[0]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(s_axi_wdata[1]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(s_axi_wdata[2]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(s_axi_wdata[3]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(s_axi_wdata[4]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(s_axi_wdata[5]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(s_axi_wdata[6]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(s_axi_wdata[7]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(s_axi_wvalid),
    .X(net22));
 sky130_fd_sc_hd__buf_4 output23 (.A(net23),
    .X(s_axi_arready));
 sky130_fd_sc_hd__buf_4 output24 (.A(net24),
    .X(s_axi_awready));
 sky130_fd_sc_hd__buf_4 output25 (.A(net25),
    .X(s_axi_bvalid));
 sky130_fd_sc_hd__buf_4 output26 (.A(net26),
    .X(s_axi_rdata[0]));
 sky130_fd_sc_hd__buf_4 output27 (.A(net27),
    .X(s_axi_rdata[1]));
 sky130_fd_sc_hd__buf_4 output28 (.A(net28),
    .X(s_axi_rdata[2]));
 sky130_fd_sc_hd__buf_4 output29 (.A(net29),
    .X(s_axi_rdata[3]));
 sky130_fd_sc_hd__buf_4 output30 (.A(net30),
    .X(s_axi_rdata[4]));
 sky130_fd_sc_hd__buf_4 output31 (.A(net31),
    .X(s_axi_rdata[5]));
 sky130_fd_sc_hd__buf_4 output32 (.A(net32),
    .X(s_axi_rdata[6]));
 sky130_fd_sc_hd__buf_4 output33 (.A(net33),
    .X(s_axi_rdata[7]));
 sky130_fd_sc_hd__buf_4 output34 (.A(net34),
    .X(s_axi_rvalid));
 sky130_fd_sc_hd__buf_4 output35 (.A(net35),
    .X(s_axi_wready));
 sky130_fd_sc_hd__buf_4 fanout36 (.A(net38),
    .X(net36));
 sky130_fd_sc_hd__buf_4 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net1),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(net1),
    .X(net40));
 sky130_fd_sc_hd__conb_1 lfsr_axi_top_41 (.LO(net41));
 assign s_axi_bresp[0] = net41;
 assign s_axi_bresp[1] = net42;
endmodule
