VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO lfsr_axi_top
  CLASS BLOCK ;
  FOREIGN lfsr_axi_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 97.940 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 105.200 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 96.340 105.200 97.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.600 -0.020 105.200 97.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.115 -0.020 20.715 97.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.310 -0.020 42.910 97.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.505 -0.020 65.105 97.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.700 -0.020 87.300 97.940 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 22.900 105.200 24.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 41.940 105.200 43.540 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 60.980 105.200 62.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 80.020 105.200 81.620 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 94.640 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 101.900 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 93.040 101.900 94.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.300 3.280 101.900 94.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.815 -0.020 17.415 97.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 -0.020 39.610 97.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 -0.020 61.805 97.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.400 -0.020 84.000 97.940 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 19.600 105.200 21.200 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 38.640 105.200 40.240 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 57.680 105.200 59.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 76.720 105.200 78.320 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END clk
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END rst_n
  PIN s_axi_araddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END s_axi_araddr[0]
  PIN s_axi_araddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END s_axi_araddr[1]
  PIN s_axi_araddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END s_axi_araddr[2]
  PIN s_axi_araddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END s_axi_araddr[3]
  PIN s_axi_arready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END s_axi_arready
  PIN s_axi_arvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END s_axi_arvalid
  PIN s_axi_awaddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END s_axi_awaddr[0]
  PIN s_axi_awaddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END s_axi_awaddr[1]
  PIN s_axi_awaddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END s_axi_awaddr[2]
  PIN s_axi_awaddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END s_axi_awaddr[3]
  PIN s_axi_awready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END s_axi_awready
  PIN s_axi_awvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END s_axi_awvalid
  PIN s_axi_bready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END s_axi_bready
  PIN s_axi_bresp[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END s_axi_bresp[0]
  PIN s_axi_bresp[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END s_axi_bresp[1]
  PIN s_axi_bvalid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END s_axi_bvalid
  PIN s_axi_rdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END s_axi_rdata[0]
  PIN s_axi_rdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END s_axi_rdata[1]
  PIN s_axi_rdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END s_axi_rdata[2]
  PIN s_axi_rdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END s_axi_rdata[3]
  PIN s_axi_rdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END s_axi_rdata[4]
  PIN s_axi_rdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END s_axi_rdata[5]
  PIN s_axi_rdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END s_axi_rdata[6]
  PIN s_axi_rdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END s_axi_rdata[7]
  PIN s_axi_rready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END s_axi_rready
  PIN s_axi_rvalid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END s_axi_rvalid
  PIN s_axi_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END s_axi_wdata[0]
  PIN s_axi_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.040 4.000 0.640 ;
    END
  END s_axi_wdata[1]
  PIN s_axi_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END s_axi_wdata[2]
  PIN s_axi_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END s_axi_wdata[3]
  PIN s_axi_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END s_axi_wdata[4]
  PIN s_axi_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END s_axi_wdata[5]
  PIN s_axi_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END s_axi_wdata[6]
  PIN s_axi_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END s_axi_wdata[7]
  PIN s_axi_wready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END s_axi_wready
  PIN s_axi_wvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END s_axi_wvalid
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 94.490 87.125 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 1.910 9.220 97.450 88.360 ;
      LAYER met2 ;
        RECT 1.930 4.280 97.420 95.725 ;
        RECT 1.930 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 97.420 4.280 ;
      LAYER met3 ;
        RECT 4.400 98.240 96.995 99.100 ;
        RECT 1.905 96.240 96.995 98.240 ;
        RECT 4.400 94.840 96.995 96.240 ;
        RECT 1.905 92.840 96.995 94.840 ;
        RECT 4.400 91.440 96.995 92.840 ;
        RECT 1.905 89.440 96.995 91.440 ;
        RECT 4.400 88.040 96.995 89.440 ;
        RECT 1.905 86.040 96.995 88.040 ;
        RECT 4.400 84.640 96.995 86.040 ;
        RECT 1.905 82.640 96.995 84.640 ;
        RECT 4.400 81.240 96.995 82.640 ;
        RECT 1.905 79.240 96.995 81.240 ;
        RECT 4.400 77.840 96.995 79.240 ;
        RECT 1.905 75.840 96.995 77.840 ;
        RECT 4.400 74.440 96.995 75.840 ;
        RECT 1.905 72.440 96.995 74.440 ;
        RECT 4.400 71.040 96.995 72.440 ;
        RECT 1.905 69.040 96.995 71.040 ;
        RECT 4.400 67.640 96.995 69.040 ;
        RECT 1.905 65.640 96.995 67.640 ;
        RECT 4.400 64.240 96.995 65.640 ;
        RECT 1.905 62.240 96.995 64.240 ;
        RECT 4.400 60.840 96.995 62.240 ;
        RECT 1.905 58.840 96.995 60.840 ;
        RECT 4.400 57.440 96.995 58.840 ;
        RECT 1.905 55.440 96.995 57.440 ;
        RECT 4.400 54.040 96.995 55.440 ;
        RECT 1.905 52.040 96.995 54.040 ;
        RECT 4.400 50.640 96.995 52.040 ;
        RECT 1.905 48.640 96.995 50.640 ;
        RECT 4.400 47.240 96.995 48.640 ;
        RECT 1.905 45.240 96.995 47.240 ;
        RECT 4.400 43.840 96.995 45.240 ;
        RECT 1.905 41.840 96.995 43.840 ;
        RECT 4.400 40.440 96.995 41.840 ;
        RECT 1.905 38.440 96.995 40.440 ;
        RECT 4.400 37.040 96.995 38.440 ;
        RECT 1.905 35.040 96.995 37.040 ;
        RECT 4.400 33.640 96.995 35.040 ;
        RECT 1.905 31.640 96.995 33.640 ;
        RECT 4.400 30.240 96.995 31.640 ;
        RECT 1.905 28.240 96.995 30.240 ;
        RECT 4.400 26.840 96.995 28.240 ;
        RECT 1.905 24.840 96.995 26.840 ;
        RECT 4.400 23.440 96.995 24.840 ;
        RECT 1.905 21.440 96.995 23.440 ;
        RECT 4.400 20.040 96.995 21.440 ;
        RECT 1.905 18.040 96.995 20.040 ;
        RECT 4.400 16.640 96.995 18.040 ;
        RECT 1.905 14.640 96.995 16.640 ;
        RECT 4.400 13.240 96.995 14.640 ;
        RECT 1.905 11.240 96.995 13.240 ;
        RECT 4.400 9.840 96.995 11.240 ;
        RECT 1.905 7.840 96.995 9.840 ;
        RECT 4.400 6.440 96.995 7.840 ;
        RECT 1.905 4.440 96.995 6.440 ;
        RECT 4.400 3.040 96.995 4.440 ;
        RECT 1.905 1.040 96.995 3.040 ;
        RECT 4.400 0.175 96.995 1.040 ;
      LAYER met4 ;
        RECT 3.975 98.340 89.865 99.105 ;
        RECT 3.975 14.455 15.415 98.340 ;
        RECT 17.815 14.455 18.715 98.340 ;
        RECT 21.115 14.455 37.610 98.340 ;
        RECT 40.010 14.455 40.910 98.340 ;
        RECT 43.310 14.455 59.805 98.340 ;
        RECT 62.205 14.455 63.105 98.340 ;
        RECT 65.505 14.455 82.000 98.340 ;
        RECT 84.400 14.455 85.300 98.340 ;
        RECT 87.700 14.455 89.865 98.340 ;
  END
END lfsr_axi_top
END LIBRARY

