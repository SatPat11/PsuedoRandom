magic
tech sky130A
magscale 1 2
timestamp 1750956226
<< checkpaint >>
rect -5008 -3936 24972 23780
<< viali >>
rect 2605 17289 2639 17323
rect 7389 17289 7423 17323
rect 7665 17289 7699 17323
rect 6745 17221 6779 17255
rect 8677 17221 8711 17255
rect 12173 17221 12207 17255
rect 14289 17221 14323 17255
rect 1409 17153 1443 17187
rect 1961 17153 1995 17187
rect 2513 17153 2547 17187
rect 2789 17153 2823 17187
rect 3065 17153 3099 17187
rect 6009 17153 6043 17187
rect 6601 17153 6635 17187
rect 6837 17153 6871 17187
rect 7021 17153 7055 17187
rect 7481 17177 7515 17211
rect 8033 17153 8067 17187
rect 11805 17153 11839 17187
rect 11989 17153 12023 17187
rect 12449 17153 12483 17187
rect 13093 17153 13127 17187
rect 1685 17085 1719 17119
rect 5365 17085 5399 17119
rect 5641 17085 5675 17119
rect 12909 17085 12943 17119
rect 13277 17085 13311 17119
rect 2145 17017 2179 17051
rect 6469 17017 6503 17051
rect 2329 16949 2363 16983
rect 2881 16949 2915 16983
rect 3617 16949 3651 16983
rect 3893 16949 3927 16983
rect 5825 16949 5859 16983
rect 8401 16949 8435 16983
rect 9137 16949 9171 16983
rect 11253 16949 11287 16983
rect 13461 16949 13495 16983
rect 13737 16949 13771 16983
rect 16313 16949 16347 16983
rect 5825 16745 5859 16779
rect 6101 16745 6135 16779
rect 7297 16745 7331 16779
rect 16037 16745 16071 16779
rect 16405 16745 16439 16779
rect 13369 16677 13403 16711
rect 13829 16677 13863 16711
rect 2053 16609 2087 16643
rect 3065 16609 3099 16643
rect 3249 16609 3283 16643
rect 4077 16609 4111 16643
rect 4169 16609 4203 16643
rect 4905 16609 4939 16643
rect 8401 16609 8435 16643
rect 8769 16609 8803 16643
rect 9873 16609 9907 16643
rect 14933 16609 14967 16643
rect 15117 16609 15151 16643
rect 15761 16609 15795 16643
rect 16497 16609 16531 16643
rect 1869 16541 1903 16575
rect 2145 16541 2179 16575
rect 3617 16541 3651 16575
rect 4721 16541 4755 16575
rect 8309 16541 8343 16575
rect 8585 16541 8619 16575
rect 9224 16541 9258 16575
rect 9321 16541 9355 16575
rect 9413 16541 9447 16575
rect 9597 16541 9631 16575
rect 11161 16541 11195 16575
rect 12081 16541 12115 16575
rect 12265 16541 12299 16575
rect 12501 16541 12535 16575
rect 16405 16541 16439 16575
rect 16681 16541 16715 16575
rect 4261 16473 4295 16507
rect 6837 16473 6871 16507
rect 7941 16473 7975 16507
rect 11529 16473 11563 16507
rect 12357 16473 12391 16507
rect 14381 16473 14415 16507
rect 15025 16473 15059 16507
rect 2605 16405 2639 16439
rect 2973 16405 3007 16439
rect 3433 16405 3467 16439
rect 4629 16405 4663 16439
rect 6561 16405 6595 16439
rect 9037 16405 9071 16439
rect 10333 16405 10367 16439
rect 11897 16405 11931 16439
rect 12641 16405 12675 16439
rect 13093 16405 13127 16439
rect 14555 16405 14589 16439
rect 16865 16405 16899 16439
rect 7113 16201 7147 16235
rect 12449 16201 12483 16235
rect 14105 16201 14139 16235
rect 15393 16201 15427 16235
rect 15577 16201 15611 16235
rect 16129 16201 16163 16235
rect 12081 16133 12115 16167
rect 1869 16065 1903 16099
rect 2789 16065 2823 16099
rect 2973 16065 3007 16099
rect 6745 16065 6779 16099
rect 8672 16065 8706 16099
rect 8769 16065 8803 16099
rect 8861 16065 8895 16099
rect 9044 16065 9078 16099
rect 9137 16065 9171 16099
rect 12725 16065 12759 16099
rect 13277 16065 13311 16099
rect 14289 16065 14323 16099
rect 15761 16065 15795 16099
rect 1593 15997 1627 16031
rect 2513 15997 2547 16031
rect 3341 15997 3375 16031
rect 6561 15997 6595 16031
rect 6653 15997 6687 16031
rect 7389 15997 7423 16031
rect 7941 15997 7975 16031
rect 11805 15997 11839 16031
rect 11989 15997 12023 16031
rect 13093 15997 13127 16031
rect 8493 15929 8527 15963
rect 9413 15929 9447 15963
rect 12541 15929 12575 15963
rect 5089 15861 5123 15895
rect 5457 15861 5491 15895
rect 5825 15861 5859 15895
rect 8217 15861 8251 15895
rect 9873 15861 9907 15895
rect 11253 15861 11287 15895
rect 13645 15861 13679 15895
rect 2237 15657 2271 15691
rect 4353 15657 4387 15691
rect 5089 15657 5123 15691
rect 7941 15657 7975 15691
rect 17233 15657 17267 15691
rect 1593 15589 1627 15623
rect 2881 15521 2915 15555
rect 6837 15521 6871 15555
rect 7205 15521 7239 15555
rect 7481 15521 7515 15555
rect 11713 15521 11747 15555
rect 1409 15453 1443 15487
rect 3249 15453 3283 15487
rect 4721 15453 4755 15487
rect 12081 15453 12115 15487
rect 17601 15453 17635 15487
rect 17785 15453 17819 15487
rect 17877 15453 17911 15487
rect 18061 15453 18095 15487
rect 18153 15453 18187 15487
rect 2605 15385 2639 15419
rect 4077 15385 4111 15419
rect 13553 15385 13587 15419
rect 8401 15317 8435 15351
rect 11529 15317 11563 15351
rect 13921 15317 13955 15351
rect 14289 15317 14323 15351
rect 14657 15317 14691 15351
rect 15025 15317 15059 15351
rect 18337 15317 18371 15351
rect 1869 15113 1903 15147
rect 8033 15113 8067 15147
rect 9321 15113 9355 15147
rect 15945 15113 15979 15147
rect 17693 15113 17727 15147
rect 5963 15045 5997 15079
rect 12265 15045 12299 15079
rect 14289 15045 14323 15079
rect 1777 14977 1811 15011
rect 2421 14977 2455 15011
rect 4997 14977 5031 15011
rect 5181 14977 5215 15011
rect 5549 14977 5583 15011
rect 6652 14977 6686 15011
rect 6745 14977 6779 15011
rect 6837 14977 6871 15011
rect 7021 14977 7055 15011
rect 7389 14977 7423 15011
rect 7757 14977 7791 15011
rect 8033 14977 8067 15011
rect 8677 14967 8711 15001
rect 8860 14980 8894 15014
rect 8953 14977 8987 15011
rect 9229 14977 9263 15011
rect 14197 14977 14231 15011
rect 14381 14977 14415 15011
rect 1685 14909 1719 14943
rect 2697 14909 2731 14943
rect 4721 14909 4755 14943
rect 7481 14909 7515 14943
rect 8217 14909 8251 14943
rect 9045 14909 9079 14943
rect 11989 14909 12023 14943
rect 15577 14909 15611 14943
rect 4169 14841 4203 14875
rect 6377 14841 6411 14875
rect 14565 14841 14599 14875
rect 2237 14773 2271 14807
rect 4629 14773 4663 14807
rect 5917 14773 5951 14807
rect 6101 14773 6135 14807
rect 8585 14773 8619 14807
rect 13737 14773 13771 14807
rect 14013 14773 14047 14807
rect 14933 14773 14967 14807
rect 15301 14773 15335 14807
rect 3065 14569 3099 14603
rect 3525 14569 3559 14603
rect 5917 14569 5951 14603
rect 7205 14569 7239 14603
rect 7573 14569 7607 14603
rect 14565 14569 14599 14603
rect 7941 14501 7975 14535
rect 8401 14501 8435 14535
rect 15025 14501 15059 14535
rect 15669 14501 15703 14535
rect 2697 14433 2731 14467
rect 4169 14433 4203 14467
rect 8677 14433 8711 14467
rect 9321 14433 9355 14467
rect 13461 14433 13495 14467
rect 16129 14433 16163 14467
rect 16221 14433 16255 14467
rect 1409 14365 1443 14399
rect 2237 14365 2271 14399
rect 6469 14365 6503 14399
rect 7205 14365 7239 14399
rect 7389 14365 7423 14399
rect 8953 14365 8987 14399
rect 10793 14365 10827 14399
rect 14105 14365 14139 14399
rect 14381 14365 14415 14399
rect 15577 14365 15611 14399
rect 4445 14297 4479 14331
rect 11529 14297 11563 14331
rect 13185 14297 13219 14331
rect 1593 14229 1627 14263
rect 1869 14229 1903 14263
rect 4077 14229 4111 14263
rect 6745 14229 6779 14263
rect 11713 14229 11747 14263
rect 13829 14229 13863 14263
rect 14197 14229 14231 14263
rect 15393 14229 15427 14263
rect 16037 14229 16071 14263
rect 1593 14025 1627 14059
rect 5733 14025 5767 14059
rect 14473 14025 14507 14059
rect 16865 14025 16899 14059
rect 4445 13957 4479 13991
rect 6101 13957 6135 13991
rect 7757 13957 7791 13991
rect 14105 13957 14139 13991
rect 1409 13889 1443 13923
rect 2789 13889 2823 13923
rect 3249 13889 3283 13923
rect 3525 13889 3559 13923
rect 4077 13889 4111 13923
rect 4170 13889 4204 13923
rect 4353 13889 4387 13923
rect 4583 13889 4617 13923
rect 9505 13889 9539 13923
rect 9874 13892 9908 13926
rect 10057 13889 10091 13923
rect 13369 13889 13403 13923
rect 2053 13821 2087 13855
rect 3341 13821 3375 13855
rect 3985 13821 4019 13855
rect 5365 13821 5399 13855
rect 9321 13821 9355 13855
rect 9689 13821 9723 13855
rect 9781 13821 9815 13855
rect 14657 13821 14691 13855
rect 14933 13821 14967 13855
rect 16405 13821 16439 13855
rect 9229 13753 9263 13787
rect 10425 13753 10459 13787
rect 2421 13685 2455 13719
rect 4721 13685 4755 13719
rect 7021 13685 7055 13719
rect 8861 13685 8895 13719
rect 11805 13685 11839 13719
rect 13737 13685 13771 13719
rect 2145 13481 2179 13515
rect 13645 13481 13679 13515
rect 14289 13481 14323 13515
rect 7849 13413 7883 13447
rect 13369 13413 13403 13447
rect 16221 13413 16255 13447
rect 2881 13345 2915 13379
rect 4537 13345 4571 13379
rect 6285 13345 6319 13379
rect 11621 13345 11655 13379
rect 14749 13345 14783 13379
rect 15393 13345 15427 13379
rect 17049 13345 17083 13379
rect 1409 13277 1443 13311
rect 1869 13277 1903 13311
rect 1961 13277 1995 13311
rect 4261 13277 4295 13311
rect 11713 13277 11747 13311
rect 11878 13277 11912 13311
rect 11989 13277 12023 13311
rect 12081 13277 12115 13311
rect 12265 13277 12299 13311
rect 15117 13277 15151 13311
rect 15300 13277 15334 13311
rect 15485 13277 15519 13311
rect 15669 13277 15703 13311
rect 16405 13277 16439 13311
rect 3617 13209 3651 13243
rect 3985 13209 4019 13243
rect 6009 13209 6043 13243
rect 11253 13209 11287 13243
rect 12725 13209 12759 13243
rect 16681 13209 16715 13243
rect 1593 13141 1627 13175
rect 1685 13141 1719 13175
rect 2513 13141 2547 13175
rect 9137 13141 9171 13175
rect 9505 13141 9539 13175
rect 12357 13141 12391 13175
rect 15761 13141 15795 13175
rect 17509 13141 17543 13175
rect 9229 12937 9263 12971
rect 9965 12937 9999 12971
rect 13921 12937 13955 12971
rect 15945 12937 15979 12971
rect 17325 12937 17359 12971
rect 5273 12869 5307 12903
rect 7941 12869 7975 12903
rect 8401 12869 8435 12903
rect 8493 12869 8527 12903
rect 10057 12869 10091 12903
rect 14289 12869 14323 12903
rect 14381 12869 14415 12903
rect 16773 12869 16807 12903
rect 17877 12869 17911 12903
rect 1501 12801 1535 12835
rect 3433 12801 3467 12835
rect 5641 12801 5675 12835
rect 5733 12801 5767 12835
rect 8304 12801 8338 12835
rect 8677 12801 8711 12835
rect 9597 12801 9631 12835
rect 14013 12801 14047 12835
rect 14106 12801 14140 12835
rect 14519 12801 14553 12835
rect 15485 12801 15519 12835
rect 16037 12801 16071 12835
rect 17233 12801 17267 12835
rect 17509 12801 17543 12835
rect 1869 12733 1903 12767
rect 3801 12733 3835 12767
rect 5549 12733 5583 12767
rect 6929 12733 6963 12767
rect 9873 12733 9907 12767
rect 11805 12733 11839 12767
rect 12173 12733 12207 12767
rect 15301 12733 15335 12767
rect 16221 12733 16255 12767
rect 17049 12733 17083 12767
rect 15117 12665 15151 12699
rect 15577 12665 15611 12699
rect 3249 12597 3283 12631
rect 6101 12597 6135 12631
rect 6653 12597 6687 12631
rect 7573 12597 7607 12631
rect 8125 12597 8159 12631
rect 10425 12597 10459 12631
rect 14657 12597 14691 12631
rect 5365 12393 5399 12427
rect 13461 12393 13495 12427
rect 17417 12393 17451 12427
rect 3617 12257 3651 12291
rect 4353 12257 4387 12291
rect 5089 12257 5123 12291
rect 8401 12257 8435 12291
rect 10793 12257 10827 12291
rect 15945 12257 15979 12291
rect 1869 12189 1903 12223
rect 2145 12189 2179 12223
rect 2329 12189 2363 12223
rect 4261 12189 4295 12223
rect 4629 12189 4663 12223
rect 4905 12189 4939 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 11069 12189 11103 12223
rect 11805 12189 11839 12223
rect 14381 12189 14415 12223
rect 15669 12189 15703 12223
rect 1593 12121 1627 12155
rect 2605 12121 2639 12155
rect 7757 12121 7791 12155
rect 10517 12121 10551 12155
rect 1961 12053 1995 12087
rect 3065 12053 3099 12087
rect 5089 12053 5123 12087
rect 5733 12053 5767 12087
rect 6469 12053 6503 12087
rect 8309 12053 8343 12087
rect 9045 12053 9079 12087
rect 10977 12053 11011 12087
rect 13921 12053 13955 12087
rect 14657 12053 14691 12087
rect 15393 12053 15427 12087
rect 6469 11849 6503 11883
rect 7941 11849 7975 11883
rect 16773 11849 16807 11883
rect 2605 11781 2639 11815
rect 3341 11781 3375 11815
rect 14105 11781 14139 11815
rect 16221 11781 16255 11815
rect 1685 11713 1719 11747
rect 1777 11713 1811 11747
rect 2416 11713 2450 11747
rect 2513 11713 2547 11747
rect 2789 11713 2823 11747
rect 3985 11713 4019 11747
rect 6561 11713 6595 11747
rect 6837 11713 6871 11747
rect 6930 11713 6964 11747
rect 7113 11713 7147 11747
rect 7573 11713 7607 11747
rect 13921 11713 13955 11747
rect 16129 11713 16163 11747
rect 16773 11713 16807 11747
rect 16957 11713 16991 11747
rect 17693 11713 17727 11747
rect 2053 11645 2087 11679
rect 4077 11645 4111 11679
rect 4169 11645 4203 11679
rect 5457 11645 5491 11679
rect 6745 11645 6779 11679
rect 7297 11645 7331 11679
rect 7481 11645 7515 11679
rect 8401 11645 8435 11679
rect 10701 11645 10735 11679
rect 13277 11645 13311 11679
rect 13461 11645 13495 11679
rect 15853 11645 15887 11679
rect 16221 11645 16255 11679
rect 16405 11645 16439 11679
rect 16497 11645 16531 11679
rect 1501 11577 1535 11611
rect 3617 11577 3651 11611
rect 1961 11509 1995 11543
rect 2237 11509 2271 11543
rect 4905 11509 4939 11543
rect 5733 11509 5767 11543
rect 6193 11509 6227 11543
rect 8861 11509 8895 11543
rect 13001 11509 13035 11543
rect 13645 11509 13679 11543
rect 17325 11509 17359 11543
rect 4353 11305 4387 11339
rect 5825 11305 5859 11339
rect 9137 11305 9171 11339
rect 11437 11305 11471 11339
rect 15209 11305 15243 11339
rect 15945 11305 15979 11339
rect 1593 11237 1627 11271
rect 4721 11237 4755 11271
rect 16957 11237 16991 11271
rect 3341 11169 3375 11203
rect 3617 11169 3651 11203
rect 7566 11169 7600 11203
rect 14473 11169 14507 11203
rect 1409 11101 1443 11135
rect 7665 11101 7699 11135
rect 7849 11101 7883 11135
rect 8125 11101 8159 11135
rect 8321 11101 8355 11135
rect 8677 11101 8711 11135
rect 12909 11101 12943 11135
rect 14197 11101 14231 11135
rect 14362 11101 14396 11135
rect 14565 11101 14599 11135
rect 14749 11101 14783 11135
rect 14933 11101 14967 11135
rect 16313 11101 16347 11135
rect 16497 11101 16531 11135
rect 16589 11101 16623 11135
rect 16715 11101 16749 11135
rect 17693 11101 17727 11135
rect 5365 11033 5399 11067
rect 7297 11033 7331 11067
rect 13553 11033 13587 11067
rect 13737 11033 13771 11067
rect 15577 11033 15611 11067
rect 17325 11033 17359 11067
rect 1869 10965 1903 10999
rect 5089 10965 5123 10999
rect 8033 10965 8067 10999
rect 1869 10761 1903 10795
rect 2881 10761 2915 10795
rect 3709 10761 3743 10795
rect 7297 10761 7331 10795
rect 10609 10761 10643 10795
rect 11253 10761 11287 10795
rect 11989 10761 12023 10795
rect 18061 10761 18095 10795
rect 2513 10693 2547 10727
rect 3617 10693 3651 10727
rect 7113 10693 7147 10727
rect 11897 10693 11931 10727
rect 14933 10693 14967 10727
rect 1409 10625 1443 10659
rect 2237 10625 2271 10659
rect 4169 10625 4203 10659
rect 6193 10625 6227 10659
rect 8585 10625 8619 10659
rect 9137 10625 9171 10659
rect 9413 10625 9447 10659
rect 9689 10625 9723 10659
rect 12817 10625 12851 10659
rect 14473 10625 14507 10659
rect 16865 10625 16899 10659
rect 17969 10625 18003 10659
rect 18337 10625 18371 10659
rect 2145 10557 2179 10591
rect 3433 10557 3467 10591
rect 4445 10557 4479 10591
rect 10241 10557 10275 10591
rect 12081 10557 12115 10591
rect 17509 10557 17543 10591
rect 18521 10557 18555 10591
rect 1593 10489 1627 10523
rect 4077 10489 4111 10523
rect 7481 10489 7515 10523
rect 8493 10489 8527 10523
rect 2237 10421 2271 10455
rect 7297 10421 7331 10455
rect 8217 10421 8251 10455
rect 11529 10421 11563 10455
rect 16037 10421 16071 10455
rect 16405 10421 16439 10455
rect 3157 10217 3191 10251
rect 3617 10217 3651 10251
rect 6285 10217 6319 10251
rect 9321 10217 9355 10251
rect 13921 10217 13955 10251
rect 4629 10149 4663 10183
rect 4721 10149 4755 10183
rect 10793 10149 10827 10183
rect 11713 10149 11747 10183
rect 4813 10081 4847 10115
rect 5917 10081 5951 10115
rect 17233 10081 17267 10115
rect 1593 10013 1627 10047
rect 1685 10013 1719 10047
rect 1961 10013 1995 10047
rect 2881 10013 2915 10047
rect 4261 10013 4295 10047
rect 7481 10013 7515 10047
rect 7677 10013 7711 10047
rect 9505 10013 9539 10047
rect 11345 10013 11379 10047
rect 11529 10013 11563 10047
rect 11713 10013 11747 10047
rect 12449 10013 12483 10047
rect 12633 10013 12667 10047
rect 13277 10013 13311 10047
rect 16405 10013 16439 10047
rect 16957 10013 16991 10047
rect 17325 10013 17359 10047
rect 17601 10013 17635 10047
rect 17969 10013 18003 10047
rect 1869 9945 1903 9979
rect 2605 9945 2639 9979
rect 5641 9945 5675 9979
rect 8309 9945 8343 9979
rect 12909 9945 12943 9979
rect 14381 9945 14415 9979
rect 16129 9945 16163 9979
rect 4077 9877 4111 9911
rect 5089 9877 5123 9911
rect 5365 9877 5399 9911
rect 5549 9877 5583 9911
rect 5733 9877 5767 9911
rect 6653 9877 6687 9911
rect 12265 9877 12299 9911
rect 8953 9673 8987 9707
rect 13829 9673 13863 9707
rect 14105 9673 14139 9707
rect 1685 9605 1719 9639
rect 3709 9605 3743 9639
rect 4813 9605 4847 9639
rect 11529 9605 11563 9639
rect 3433 9537 3467 9571
rect 5089 9537 5123 9571
rect 10776 9537 10810 9571
rect 10925 9537 10959 9571
rect 11069 9537 11103 9571
rect 11161 9537 11195 9571
rect 11345 9537 11379 9571
rect 13645 9537 13679 9571
rect 14289 9537 14323 9571
rect 14565 9537 14599 9571
rect 14933 9537 14967 9571
rect 16737 9537 16771 9571
rect 17141 9537 17175 9571
rect 17693 9537 17727 9571
rect 17785 9537 17819 9571
rect 1409 9469 1443 9503
rect 7205 9469 7239 9503
rect 7481 9469 7515 9503
rect 10241 9469 10275 9503
rect 13553 9469 13587 9503
rect 14105 9469 14139 9503
rect 15117 9469 15151 9503
rect 15393 9469 15427 9503
rect 16841 9469 16875 9503
rect 17325 9469 17359 9503
rect 18061 9469 18095 9503
rect 18337 9469 18371 9503
rect 4169 9401 4203 9435
rect 9505 9401 9539 9435
rect 9873 9401 9907 9435
rect 15761 9401 15795 9435
rect 5549 9333 5583 9367
rect 10609 9333 10643 9367
rect 13289 9333 13323 9367
rect 16221 9333 16255 9367
rect 17509 9333 17543 9367
rect 17969 9333 18003 9367
rect 2329 9129 2363 9163
rect 2513 9129 2547 9163
rect 2881 9129 2915 9163
rect 5273 9129 5307 9163
rect 6193 9129 6227 9163
rect 10333 9129 10367 9163
rect 15209 9129 15243 9163
rect 15761 9129 15795 9163
rect 10977 9061 11011 9095
rect 11161 9061 11195 9095
rect 4629 8993 4663 9027
rect 5733 8993 5767 9027
rect 5825 8993 5859 9027
rect 8493 8993 8527 9027
rect 13001 8993 13035 9027
rect 13369 8993 13403 9027
rect 16037 8993 16071 9027
rect 16497 8993 16531 9027
rect 18245 8993 18279 9027
rect 1409 8925 1443 8959
rect 2421 8925 2455 8959
rect 4353 8925 4387 8959
rect 6009 8925 6043 8959
rect 8769 8925 8803 8959
rect 9229 8925 9263 8959
rect 9597 8925 9631 8959
rect 9965 8925 9999 8959
rect 10333 8925 10367 8959
rect 12541 8925 12575 8959
rect 12909 8925 12943 8959
rect 14105 8925 14139 8959
rect 16405 8925 16439 8959
rect 6285 8857 6319 8891
rect 13461 8857 13495 8891
rect 13737 8857 13771 8891
rect 16773 8857 16807 8891
rect 3985 8789 4019 8823
rect 4445 8789 4479 8823
rect 7021 8789 7055 8823
rect 13277 8789 13311 8823
rect 14289 8789 14323 8823
rect 14657 8789 14691 8823
rect 16221 8789 16255 8823
rect 8953 8585 8987 8619
rect 13737 8585 13771 8619
rect 14013 8585 14047 8619
rect 15117 8585 15151 8619
rect 15853 8585 15887 8619
rect 16865 8585 16899 8619
rect 18429 8585 18463 8619
rect 3801 8517 3835 8551
rect 8125 8517 8159 8551
rect 11529 8517 11563 8551
rect 15761 8517 15795 8551
rect 18153 8517 18187 8551
rect 1593 8449 1627 8483
rect 2145 8449 2179 8483
rect 5825 8449 5859 8483
rect 6377 8449 6411 8483
rect 9321 8449 9355 8483
rect 11345 8449 11379 8483
rect 17049 8449 17083 8483
rect 17785 8449 17819 8483
rect 17878 8449 17912 8483
rect 18061 8449 18095 8483
rect 18291 8449 18325 8483
rect 1685 8381 1719 8415
rect 1777 8381 1811 8415
rect 5549 8381 5583 8415
rect 9597 8381 9631 8415
rect 13001 8381 13035 8415
rect 13369 8381 13403 8415
rect 16037 8381 16071 8415
rect 16405 8381 16439 8415
rect 17141 8381 17175 8415
rect 17325 8381 17359 8415
rect 17509 8381 17543 8415
rect 15393 8313 15427 8347
rect 2421 8245 2455 8279
rect 14749 8245 14783 8279
rect 2697 8041 2731 8075
rect 3157 8041 3191 8075
rect 6377 8041 6411 8075
rect 9873 8041 9907 8075
rect 13921 8041 13955 8075
rect 15669 8041 15703 8075
rect 16313 8041 16347 8075
rect 9137 7973 9171 8007
rect 15025 7973 15059 8007
rect 16773 7973 16807 8007
rect 17693 7973 17727 8007
rect 1593 7905 1627 7939
rect 8677 7905 8711 7939
rect 9505 7905 9539 7939
rect 10701 7905 10735 7939
rect 14841 7905 14875 7939
rect 1869 7837 1903 7871
rect 2421 7837 2455 7871
rect 4077 7837 4111 7871
rect 4445 7837 4479 7871
rect 4813 7837 4847 7871
rect 5089 7837 5123 7871
rect 5549 7837 5583 7871
rect 9321 7837 9355 7871
rect 10977 7837 11011 7871
rect 15025 7837 15059 7871
rect 15669 7837 15703 7871
rect 16037 7837 16071 7871
rect 17325 7837 17359 7871
rect 18245 7837 18279 7871
rect 2145 7769 2179 7803
rect 4997 7769 5031 7803
rect 10057 7769 10091 7803
rect 15393 7769 15427 7803
rect 5917 7701 5951 7735
rect 9689 7701 9723 7735
rect 9873 7701 9907 7735
rect 10333 7701 10367 7735
rect 11345 7701 11379 7735
rect 11621 7701 11655 7735
rect 13461 7701 13495 7735
rect 14289 7701 14323 7735
rect 14749 7701 14783 7735
rect 15853 7701 15887 7735
rect 17141 7701 17175 7735
rect 18061 7701 18095 7735
rect 9229 7497 9263 7531
rect 10793 7497 10827 7531
rect 14381 7497 14415 7531
rect 14749 7497 14783 7531
rect 17141 7497 17175 7531
rect 17509 7497 17543 7531
rect 3525 7429 3559 7463
rect 4077 7429 4111 7463
rect 9597 7429 9631 7463
rect 15393 7429 15427 7463
rect 16497 7429 16531 7463
rect 1869 7361 1903 7395
rect 9965 7361 9999 7395
rect 10333 7361 10367 7395
rect 10609 7385 10643 7419
rect 11161 7361 11195 7395
rect 12173 7361 12207 7395
rect 14289 7361 14323 7395
rect 17049 7361 17083 7395
rect 18153 7361 18187 7395
rect 18337 7361 18371 7395
rect 1593 7293 1627 7327
rect 2053 7293 2087 7327
rect 3812 7293 3846 7327
rect 10517 7293 10551 7327
rect 14105 7293 14139 7327
rect 16037 7293 16071 7327
rect 16957 7293 16991 7327
rect 17693 7293 17727 7327
rect 17877 7293 17911 7327
rect 17969 7293 18003 7327
rect 18061 7293 18095 7327
rect 5457 7225 5491 7259
rect 10057 7225 10091 7259
rect 13645 7157 13679 7191
rect 15761 7157 15795 7191
rect 2145 6953 2179 6987
rect 7125 6953 7159 6987
rect 9873 6953 9907 6987
rect 11909 6953 11943 6987
rect 14289 6953 14323 6987
rect 16681 6953 16715 6987
rect 2605 6885 2639 6919
rect 10425 6885 10459 6919
rect 12725 6885 12759 6919
rect 17877 6885 17911 6919
rect 4445 6817 4479 6851
rect 8401 6817 8435 6851
rect 12173 6817 12207 6851
rect 1869 6749 1903 6783
rect 1961 6749 1995 6783
rect 2789 6749 2823 6783
rect 4353 6749 4387 6783
rect 7389 6749 7423 6783
rect 8309 6749 8343 6783
rect 8585 6749 8619 6783
rect 12449 6749 12483 6783
rect 12909 6749 12943 6783
rect 13093 6749 13127 6783
rect 13369 6749 13403 6783
rect 17417 6749 17451 6783
rect 17785 6749 17819 6783
rect 18337 6749 18371 6783
rect 2145 6681 2179 6715
rect 3525 6681 3559 6715
rect 3801 6681 3835 6715
rect 4077 6681 4111 6715
rect 5365 6681 5399 6715
rect 12265 6681 12299 6715
rect 12633 6681 12667 6715
rect 13737 6681 13771 6715
rect 1685 6613 1719 6647
rect 2973 6613 3007 6647
rect 3433 6613 3467 6647
rect 8769 6613 8803 6647
rect 16957 6613 16991 6647
rect 3249 6409 3283 6443
rect 5273 6409 5307 6443
rect 6653 6409 6687 6443
rect 6745 6409 6779 6443
rect 7113 6409 7147 6443
rect 9689 6409 9723 6443
rect 12265 6409 12299 6443
rect 13553 6409 13587 6443
rect 17049 6409 17083 6443
rect 17509 6409 17543 6443
rect 17877 6409 17911 6443
rect 2421 6341 2455 6375
rect 5549 6341 5583 6375
rect 5641 6341 5675 6375
rect 9137 6341 9171 6375
rect 9505 6341 9539 6375
rect 10057 6341 10091 6375
rect 12909 6341 12943 6375
rect 1869 6273 1903 6307
rect 2881 6273 2915 6307
rect 5385 6273 5419 6307
rect 5738 6273 5772 6307
rect 9413 6273 9447 6307
rect 10425 6273 10459 6307
rect 12449 6273 12483 6307
rect 12541 6273 12575 6307
rect 13093 6273 13127 6307
rect 13277 6273 13311 6307
rect 1593 6205 1627 6239
rect 2697 6205 2731 6239
rect 2789 6205 2823 6239
rect 4813 6205 4847 6239
rect 6561 6205 6595 6239
rect 12817 6205 12851 6239
rect 3709 6137 3743 6171
rect 4169 6137 4203 6171
rect 5917 6137 5951 6171
rect 7665 6137 7699 6171
rect 11989 6137 12023 6171
rect 4537 6069 4571 6103
rect 7389 6069 7423 6103
rect 12725 6069 12759 6103
rect 18245 6069 18279 6103
rect 2145 5865 2179 5899
rect 2605 5865 2639 5899
rect 3985 5865 4019 5899
rect 5365 5865 5399 5899
rect 6285 5865 6319 5899
rect 7757 5865 7791 5899
rect 14197 5865 14231 5899
rect 17601 5865 17635 5899
rect 18061 5865 18095 5899
rect 7113 5797 7147 5831
rect 2237 5729 2271 5763
rect 2973 5729 3007 5763
rect 6469 5729 6503 5763
rect 12909 5729 12943 5763
rect 15945 5729 15979 5763
rect 18429 5729 18463 5763
rect 1869 5661 1903 5695
rect 1961 5661 1995 5695
rect 2053 5661 2087 5695
rect 5917 5661 5951 5695
rect 6101 5661 6135 5695
rect 8125 5661 8159 5695
rect 1593 5593 1627 5627
rect 3617 5593 3651 5627
rect 6653 5593 6687 5627
rect 8321 5593 8355 5627
rect 9413 5593 9447 5627
rect 15669 5593 15703 5627
rect 5733 5525 5767 5559
rect 6745 5525 6779 5559
rect 7481 5525 7515 5559
rect 12541 5525 12575 5559
rect 2329 5321 2363 5355
rect 10057 5321 10091 5355
rect 18153 5321 18187 5355
rect 9505 5253 9539 5287
rect 1869 5185 1903 5219
rect 2697 5185 2731 5219
rect 2973 5185 3007 5219
rect 6561 5185 6595 5219
rect 7389 5185 7423 5219
rect 9781 5185 9815 5219
rect 10241 5185 10275 5219
rect 18337 5185 18371 5219
rect 18429 5185 18463 5219
rect 1593 5117 1627 5151
rect 2789 5117 2823 5151
rect 3249 5117 3283 5151
rect 3525 5117 3559 5151
rect 5457 5117 5491 5151
rect 8033 5117 8067 5151
rect 17785 5117 17819 5151
rect 18153 5117 18187 5151
rect 4997 4981 5031 5015
rect 7757 4981 7791 5015
rect 2145 4777 2179 4811
rect 2605 4777 2639 4811
rect 3157 4777 3191 4811
rect 14197 4777 14231 4811
rect 14657 4777 14691 4811
rect 3433 4709 3467 4743
rect 4629 4709 4663 4743
rect 6101 4709 6135 4743
rect 17049 4709 17083 4743
rect 4169 4641 4203 4675
rect 5273 4641 5307 4675
rect 8769 4641 8803 4675
rect 13921 4641 13955 4675
rect 16865 4641 16899 4675
rect 1869 4573 1903 4607
rect 4261 4573 4295 4607
rect 4997 4573 5031 4607
rect 7573 4573 7607 4607
rect 8401 4573 8435 4607
rect 14289 4573 14323 4607
rect 17233 4573 17267 4607
rect 18061 4573 18095 4607
rect 1593 4505 1627 4539
rect 17877 4505 17911 4539
rect 4445 4437 4479 4471
rect 5089 4437 5123 4471
rect 5641 4437 5675 4471
rect 8008 4437 8042 4471
rect 1961 4233 1995 4267
rect 5365 4165 5399 4199
rect 2697 4097 2731 4131
rect 2973 4097 3007 4131
rect 4905 4097 4939 4131
rect 5733 4097 5767 4131
rect 6193 4097 6227 4131
rect 11069 4097 11103 4131
rect 15301 4097 15335 4131
rect 15577 4097 15611 4131
rect 17049 4097 17083 4131
rect 18521 4097 18555 4131
rect 2513 4029 2547 4063
rect 4445 4029 4479 4063
rect 4807 4029 4841 4063
rect 10793 4029 10827 4063
rect 12909 4029 12943 4063
rect 14657 4029 14691 4063
rect 14933 4029 14967 4063
rect 16681 4029 16715 4063
rect 2881 3961 2915 3995
rect 9321 3961 9355 3995
rect 12817 3893 12851 3927
rect 16405 3893 16439 3927
rect 2973 3689 3007 3723
rect 4905 3689 4939 3723
rect 6469 3689 6503 3723
rect 9873 3689 9907 3723
rect 13645 3689 13679 3723
rect 15209 3689 15243 3723
rect 15485 3689 15519 3723
rect 2697 3621 2731 3655
rect 9597 3621 9631 3655
rect 14657 3621 14691 3655
rect 1593 3553 1627 3587
rect 3617 3553 3651 3587
rect 4169 3553 4203 3587
rect 12817 3553 12851 3587
rect 14289 3553 14323 3587
rect 14933 3553 14967 3587
rect 16037 3553 16071 3587
rect 16313 3553 16347 3587
rect 18061 3553 18095 3587
rect 1869 3485 1903 3519
rect 2513 3485 2547 3519
rect 4353 3485 4387 3519
rect 4537 3485 4571 3519
rect 5365 3485 5399 3519
rect 5548 3485 5582 3519
rect 5641 3485 5675 3519
rect 5733 3485 5767 3519
rect 5917 3485 5951 3519
rect 8033 3485 8067 3519
rect 13093 3485 13127 3519
rect 13277 3485 13311 3519
rect 13466 3485 13500 3519
rect 14381 3485 14415 3519
rect 16681 3485 16715 3519
rect 6101 3417 6135 3451
rect 13369 3417 13403 3451
rect 15853 3417 15887 3451
rect 2145 3349 2179 3383
rect 3985 3349 4019 3383
rect 7849 3349 7883 3383
rect 8493 3349 8527 3383
rect 9137 3349 9171 3383
rect 12265 3349 12299 3383
rect 15945 3349 15979 3383
rect 1961 3145 1995 3179
rect 4261 3145 4295 3179
rect 4629 3145 4663 3179
rect 5273 3145 5307 3179
rect 5641 3145 5675 3179
rect 7481 3145 7515 3179
rect 10149 3145 10183 3179
rect 10333 3145 10367 3179
rect 12541 3145 12575 3179
rect 16865 3145 16899 3179
rect 17785 3145 17819 3179
rect 15669 3077 15703 3111
rect 16129 3077 16163 3111
rect 1869 3009 1903 3043
rect 2145 3009 2179 3043
rect 2605 3009 2639 3043
rect 2789 3009 2823 3043
rect 7849 3009 7883 3043
rect 8125 3009 8159 3043
rect 8677 3009 8711 3043
rect 8953 3009 8987 3043
rect 10517 3009 10551 3043
rect 10609 3009 10643 3043
rect 10701 3009 10735 3043
rect 10793 3009 10827 3043
rect 10977 3009 11011 3043
rect 12173 3009 12207 3043
rect 12357 3009 12391 3043
rect 17325 3009 17359 3043
rect 18245 3009 18279 3043
rect 1593 2941 1627 2975
rect 3065 2941 3099 2975
rect 3525 2941 3559 2975
rect 7573 2941 7607 2975
rect 9413 2941 9447 2975
rect 9781 2941 9815 2975
rect 11897 2941 11931 2975
rect 12909 2941 12943 2975
rect 13277 2941 13311 2975
rect 14657 2941 14691 2975
rect 17969 2941 18003 2975
rect 18153 2941 18187 2975
rect 2421 2873 2455 2907
rect 11253 2805 11287 2839
rect 15301 2805 15335 2839
rect 2421 2601 2455 2635
rect 4445 2601 4479 2635
rect 7297 2601 7331 2635
rect 7481 2601 7515 2635
rect 8493 2601 8527 2635
rect 10609 2601 10643 2635
rect 11069 2601 11103 2635
rect 13553 2601 13587 2635
rect 17325 2601 17359 2635
rect 17785 2601 17819 2635
rect 2145 2533 2179 2567
rect 8769 2533 8803 2567
rect 14565 2533 14599 2567
rect 15393 2533 15427 2567
rect 4077 2465 4111 2499
rect 5917 2465 5951 2499
rect 6193 2465 6227 2499
rect 7849 2465 7883 2499
rect 8033 2465 8067 2499
rect 11805 2465 11839 2499
rect 1869 2397 1903 2431
rect 1961 2397 1995 2431
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 6653 2397 6687 2431
rect 7665 2397 7699 2431
rect 8585 2397 8619 2431
rect 9137 2397 9171 2431
rect 9781 2397 9815 2431
rect 10425 2397 10459 2431
rect 11253 2397 11287 2431
rect 14289 2397 14323 2431
rect 14841 2397 14875 2431
rect 14933 2397 14967 2431
rect 15117 2397 15151 2431
rect 15209 2397 15243 2431
rect 1593 2329 1627 2363
rect 3249 2329 3283 2363
rect 12081 2329 12115 2363
rect 15761 2329 15795 2363
rect 7021 2261 7055 2295
rect 8125 2261 8159 2295
rect 9321 2261 9355 2295
rect 9965 2261 9999 2295
rect 14105 2261 14139 2295
<< metal1 >>
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 13814 17660 13820 17672
rect 6236 17632 13820 17660
rect 6236 17620 6242 17632
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 7374 17552 7380 17604
rect 7432 17592 7438 17604
rect 18966 17592 18972 17604
rect 7432 17564 18972 17592
rect 7432 17552 7438 17564
rect 18966 17552 18972 17564
rect 19024 17552 19030 17604
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 13078 17524 13084 17536
rect 6052 17496 13084 17524
rect 6052 17484 6058 17496
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 1104 17434 18860 17456
rect 1104 17382 3829 17434
rect 3881 17382 3893 17434
rect 3945 17382 3957 17434
rect 4009 17382 4021 17434
rect 4073 17382 4085 17434
rect 4137 17382 8268 17434
rect 8320 17382 8332 17434
rect 8384 17382 8396 17434
rect 8448 17382 8460 17434
rect 8512 17382 8524 17434
rect 8576 17382 12707 17434
rect 12759 17382 12771 17434
rect 12823 17382 12835 17434
rect 12887 17382 12899 17434
rect 12951 17382 12963 17434
rect 13015 17382 17146 17434
rect 17198 17382 17210 17434
rect 17262 17382 17274 17434
rect 17326 17382 17338 17434
rect 17390 17382 17402 17434
rect 17454 17382 18860 17434
rect 1104 17360 18860 17382
rect 2593 17323 2651 17329
rect 2593 17289 2605 17323
rect 2639 17320 2651 17323
rect 3694 17320 3700 17332
rect 2639 17292 3700 17320
rect 2639 17289 2651 17292
rect 2593 17283 2651 17289
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 6822 17320 6828 17332
rect 6748 17292 6828 17320
rect 2866 17252 2872 17264
rect 1964 17224 2872 17252
rect 1397 17187 1455 17193
rect 1397 17153 1409 17187
rect 1443 17184 1455 17187
rect 1486 17184 1492 17196
rect 1443 17156 1492 17184
rect 1443 17153 1455 17156
rect 1397 17147 1455 17153
rect 1486 17144 1492 17156
rect 1544 17144 1550 17196
rect 1964 17193 1992 17224
rect 2866 17212 2872 17224
rect 2924 17212 2930 17264
rect 2958 17212 2964 17264
rect 3016 17252 3022 17264
rect 3602 17252 3608 17264
rect 3016 17224 3608 17252
rect 3016 17212 3022 17224
rect 3602 17212 3608 17224
rect 3660 17212 3666 17264
rect 4338 17212 4344 17264
rect 4396 17212 4402 17264
rect 6748 17261 6776 17292
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 7374 17320 7380 17332
rect 6932 17292 7380 17320
rect 6733 17255 6791 17261
rect 6733 17221 6745 17255
rect 6779 17221 6791 17255
rect 6733 17215 6791 17221
rect 1949 17187 2007 17193
rect 1949 17153 1961 17187
rect 1995 17153 2007 17187
rect 1949 17147 2007 17153
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17184 2559 17187
rect 2777 17187 2835 17193
rect 2547 17156 2728 17184
rect 2547 17153 2559 17156
rect 2501 17147 2559 17153
rect 2700 17128 2728 17156
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 2976 17184 3004 17212
rect 2823 17156 3004 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6546 17144 6552 17196
rect 6604 17193 6610 17196
rect 6604 17187 6647 17193
rect 6635 17153 6647 17187
rect 6604 17147 6647 17153
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 6932 17184 6960 17292
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17320 7711 17323
rect 9214 17320 9220 17332
rect 7699 17292 9220 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 16942 17320 16948 17332
rect 9324 17292 16948 17320
rect 7469 17211 7527 17217
rect 7558 17212 7564 17264
rect 7616 17252 7622 17264
rect 8665 17255 8723 17261
rect 8665 17252 8677 17255
rect 7616 17224 8677 17252
rect 7616 17212 7622 17224
rect 8665 17221 8677 17224
rect 8711 17252 8723 17255
rect 9324 17252 9352 17292
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 8711 17224 9352 17252
rect 8711 17221 8723 17224
rect 8665 17215 8723 17221
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 9456 17224 12020 17252
rect 9456 17212 9462 17224
rect 7009 17188 7067 17193
rect 6871 17156 6960 17184
rect 7003 17187 7067 17188
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 7003 17153 7021 17187
rect 7055 17153 7067 17187
rect 7003 17147 7067 17153
rect 6604 17144 6610 17147
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17085 1731 17119
rect 1673 17079 1731 17085
rect 1688 17048 1716 17079
rect 2682 17076 2688 17128
rect 2740 17116 2746 17128
rect 3510 17116 3516 17128
rect 2740 17088 3516 17116
rect 2740 17076 2746 17088
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 5350 17076 5356 17128
rect 5408 17076 5414 17128
rect 5626 17076 5632 17128
rect 5684 17076 5690 17128
rect 7003 17116 7031 17147
rect 7190 17144 7196 17196
rect 7248 17184 7254 17196
rect 7469 17184 7481 17211
rect 7248 17177 7481 17184
rect 7515 17177 7527 17211
rect 7248 17171 7527 17177
rect 7248 17156 7512 17171
rect 7248 17144 7254 17156
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7708 17156 8033 17184
rect 7708 17144 7714 17156
rect 8021 17153 8033 17156
rect 8067 17184 8079 17187
rect 9766 17184 9772 17196
rect 8067 17156 9772 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 11790 17144 11796 17196
rect 11848 17144 11854 17196
rect 11992 17193 12020 17224
rect 12158 17212 12164 17264
rect 12216 17212 12222 17264
rect 12526 17212 12532 17264
rect 12584 17252 12590 17264
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 12584 17224 14289 17252
rect 12584 17212 12590 17224
rect 14277 17221 14289 17224
rect 14323 17252 14335 17255
rect 15194 17252 15200 17264
rect 14323 17224 15200 17252
rect 14323 17221 14335 17224
rect 14277 17215 14335 17221
rect 15194 17212 15200 17224
rect 15252 17212 15258 17264
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17184 12035 17187
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12023 17156 12449 17184
rect 12023 17153 12035 17156
rect 11977 17147 12035 17153
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17184 13139 17187
rect 13630 17184 13636 17196
rect 13127 17156 13636 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 8386 17116 8392 17128
rect 7003 17088 8392 17116
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 8754 17076 8760 17128
rect 8812 17116 8818 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 8812 17088 12909 17116
rect 8812 17076 8818 17088
rect 12897 17085 12909 17088
rect 12943 17116 12955 17119
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 12943 17088 13277 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 13265 17085 13277 17088
rect 13311 17116 13323 17119
rect 16022 17116 16028 17128
rect 13311 17088 16028 17116
rect 13311 17085 13323 17088
rect 13265 17079 13323 17085
rect 16022 17076 16028 17088
rect 16080 17076 16086 17128
rect 1946 17048 1952 17060
rect 1688 17020 1952 17048
rect 1946 17008 1952 17020
rect 2004 17008 2010 17060
rect 2133 17051 2191 17057
rect 2133 17017 2145 17051
rect 2179 17048 2191 17051
rect 5994 17048 6000 17060
rect 2179 17020 4384 17048
rect 2179 17017 2191 17020
rect 2133 17011 2191 17017
rect 2317 16983 2375 16989
rect 2317 16949 2329 16983
rect 2363 16980 2375 16983
rect 2682 16980 2688 16992
rect 2363 16952 2688 16980
rect 2363 16949 2375 16952
rect 2317 16943 2375 16949
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 2869 16983 2927 16989
rect 2869 16949 2881 16983
rect 2915 16980 2927 16983
rect 3050 16980 3056 16992
rect 2915 16952 3056 16980
rect 2915 16949 2927 16952
rect 2869 16943 2927 16949
rect 3050 16940 3056 16952
rect 3108 16940 3114 16992
rect 3605 16983 3663 16989
rect 3605 16949 3617 16983
rect 3651 16980 3663 16983
rect 3786 16980 3792 16992
rect 3651 16952 3792 16980
rect 3651 16949 3663 16952
rect 3605 16943 3663 16949
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 3878 16940 3884 16992
rect 3936 16940 3942 16992
rect 4356 16980 4384 17020
rect 5552 17020 6000 17048
rect 5552 16980 5580 17020
rect 5994 17008 6000 17020
rect 6052 17008 6058 17060
rect 6457 17051 6515 17057
rect 6457 17017 6469 17051
rect 6503 17048 6515 17051
rect 11146 17048 11152 17060
rect 6503 17020 11152 17048
rect 6503 17017 6515 17020
rect 6457 17011 6515 17017
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 4356 16952 5580 16980
rect 5813 16983 5871 16989
rect 5813 16949 5825 16983
rect 5859 16980 5871 16983
rect 5902 16980 5908 16992
rect 5859 16952 5908 16980
rect 5859 16949 5871 16952
rect 5813 16943 5871 16949
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 6546 16940 6552 16992
rect 6604 16980 6610 16992
rect 7098 16980 7104 16992
rect 6604 16952 7104 16980
rect 6604 16940 6610 16952
rect 7098 16940 7104 16952
rect 7156 16980 7162 16992
rect 7374 16980 7380 16992
rect 7156 16952 7380 16980
rect 7156 16940 7162 16952
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 8386 16940 8392 16992
rect 8444 16940 8450 16992
rect 8846 16940 8852 16992
rect 8904 16980 8910 16992
rect 9122 16980 9128 16992
rect 8904 16952 9128 16980
rect 8904 16940 8910 16952
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 11241 16983 11299 16989
rect 11241 16980 11253 16983
rect 10836 16952 11253 16980
rect 10836 16940 10842 16952
rect 11241 16949 11253 16952
rect 11287 16980 11299 16983
rect 11790 16980 11796 16992
rect 11287 16952 11796 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 13446 16940 13452 16992
rect 13504 16940 13510 16992
rect 13630 16940 13636 16992
rect 13688 16980 13694 16992
rect 13725 16983 13783 16989
rect 13725 16980 13737 16983
rect 13688 16952 13737 16980
rect 13688 16940 13694 16952
rect 13725 16949 13737 16952
rect 13771 16949 13783 16983
rect 13725 16943 13783 16949
rect 16298 16940 16304 16992
rect 16356 16940 16362 16992
rect 1104 16890 18860 16912
rect 1104 16838 3169 16890
rect 3221 16838 3233 16890
rect 3285 16838 3297 16890
rect 3349 16838 3361 16890
rect 3413 16838 3425 16890
rect 3477 16838 7608 16890
rect 7660 16838 7672 16890
rect 7724 16838 7736 16890
rect 7788 16838 7800 16890
rect 7852 16838 7864 16890
rect 7916 16838 12047 16890
rect 12099 16838 12111 16890
rect 12163 16838 12175 16890
rect 12227 16838 12239 16890
rect 12291 16838 12303 16890
rect 12355 16838 16486 16890
rect 16538 16838 16550 16890
rect 16602 16838 16614 16890
rect 16666 16838 16678 16890
rect 16730 16838 16742 16890
rect 16794 16838 18860 16890
rect 1104 16816 18860 16838
rect 4430 16736 4436 16788
rect 4488 16776 4494 16788
rect 4488 16748 4844 16776
rect 4488 16736 4494 16748
rect 3786 16708 3792 16720
rect 3068 16680 3792 16708
rect 2038 16600 2044 16652
rect 2096 16600 2102 16652
rect 2958 16640 2964 16652
rect 2148 16612 2964 16640
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 1946 16572 1952 16584
rect 1903 16544 1952 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 2148 16581 2176 16612
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3068 16649 3096 16680
rect 3786 16668 3792 16680
rect 3844 16708 3850 16720
rect 4338 16708 4344 16720
rect 3844 16680 4344 16708
rect 3844 16668 3850 16680
rect 4338 16668 4344 16680
rect 4396 16668 4402 16720
rect 4816 16708 4844 16748
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 5810 16776 5816 16788
rect 5592 16748 5816 16776
rect 5592 16736 5598 16748
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 5994 16736 6000 16788
rect 6052 16776 6058 16788
rect 6089 16779 6147 16785
rect 6089 16776 6101 16779
rect 6052 16748 6101 16776
rect 6052 16736 6058 16748
rect 6089 16745 6101 16748
rect 6135 16745 6147 16779
rect 6089 16739 6147 16745
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7282 16776 7288 16788
rect 6972 16748 7288 16776
rect 6972 16736 6978 16748
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 11238 16776 11244 16788
rect 9048 16748 11244 16776
rect 4816 16680 4936 16708
rect 3053 16643 3111 16649
rect 3053 16609 3065 16643
rect 3099 16609 3111 16643
rect 3053 16603 3111 16609
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 3292 16612 4077 16640
rect 3292 16600 3298 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4246 16640 4252 16652
rect 4203 16612 4252 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 2133 16535 2191 16541
rect 2774 16532 2780 16584
rect 2832 16572 2838 16584
rect 3605 16575 3663 16581
rect 3605 16572 3617 16575
rect 2832 16544 3617 16572
rect 2832 16532 2838 16544
rect 3605 16541 3617 16544
rect 3651 16541 3663 16575
rect 4080 16572 4108 16603
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 4908 16649 4936 16680
rect 4893 16643 4951 16649
rect 4356 16612 4844 16640
rect 4356 16572 4384 16612
rect 4080 16544 4384 16572
rect 3605 16535 3663 16541
rect 4706 16532 4712 16584
rect 4764 16532 4770 16584
rect 4816 16572 4844 16612
rect 4893 16609 4905 16643
rect 4939 16609 4951 16643
rect 4893 16603 4951 16609
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 5592 16612 8401 16640
rect 5592 16600 5598 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 8389 16603 8447 16609
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 8757 16643 8815 16649
rect 8757 16640 8769 16643
rect 8536 16612 8769 16640
rect 8536 16600 8542 16612
rect 8757 16609 8769 16612
rect 8803 16640 8815 16643
rect 8938 16640 8944 16652
rect 8803 16612 8944 16640
rect 8803 16609 8815 16612
rect 8757 16603 8815 16609
rect 8938 16600 8944 16612
rect 8996 16640 9002 16652
rect 9048 16640 9076 16748
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 12124 16748 12756 16776
rect 12124 16736 12130 16748
rect 9490 16668 9496 16720
rect 9548 16668 9554 16720
rect 11514 16668 11520 16720
rect 11572 16708 11578 16720
rect 12250 16708 12256 16720
rect 11572 16680 12256 16708
rect 11572 16668 11578 16680
rect 12250 16668 12256 16680
rect 12308 16668 12314 16720
rect 12728 16708 12756 16748
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 16356 16748 16405 16776
rect 16356 16736 16362 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 13357 16711 13415 16717
rect 13357 16708 13369 16711
rect 12728 16680 13369 16708
rect 13357 16677 13369 16680
rect 13403 16677 13415 16711
rect 13357 16671 13415 16677
rect 8996 16612 9076 16640
rect 8996 16600 9002 16612
rect 9122 16600 9128 16652
rect 9180 16640 9186 16652
rect 9508 16640 9536 16668
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9180 16612 9444 16640
rect 9508 16612 9873 16640
rect 9180 16600 9186 16612
rect 6638 16572 6644 16584
rect 4816 16544 6644 16572
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 8297 16575 8355 16581
rect 8297 16541 8309 16575
rect 8343 16572 8355 16575
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 8343 16544 8585 16572
rect 8343 16541 8355 16544
rect 8297 16535 8355 16541
rect 8573 16541 8585 16544
rect 8619 16572 8631 16575
rect 8662 16572 8668 16584
rect 8619 16544 8668 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8662 16532 8668 16544
rect 8720 16572 8726 16584
rect 9212 16575 9270 16581
rect 9212 16572 9224 16575
rect 8720 16544 9224 16572
rect 8720 16532 8726 16544
rect 9212 16541 9224 16544
rect 9258 16541 9270 16575
rect 9212 16535 9270 16541
rect 2222 16464 2228 16516
rect 2280 16504 2286 16516
rect 4249 16507 4307 16513
rect 2280 16476 3464 16504
rect 2280 16464 2286 16476
rect 1854 16396 1860 16448
rect 1912 16436 1918 16448
rect 2593 16439 2651 16445
rect 2593 16436 2605 16439
rect 1912 16408 2605 16436
rect 1912 16396 1918 16408
rect 2593 16405 2605 16408
rect 2639 16405 2651 16439
rect 2593 16399 2651 16405
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3436 16445 3464 16476
rect 4249 16473 4261 16507
rect 4295 16504 4307 16507
rect 4295 16476 4936 16504
rect 4295 16473 4307 16476
rect 4249 16467 4307 16473
rect 2961 16439 3019 16445
rect 2961 16436 2973 16439
rect 2832 16408 2973 16436
rect 2832 16396 2838 16408
rect 2961 16405 2973 16408
rect 3007 16405 3019 16439
rect 2961 16399 3019 16405
rect 3421 16439 3479 16445
rect 3421 16405 3433 16439
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 4614 16396 4620 16448
rect 4672 16396 4678 16448
rect 4908 16436 4936 16476
rect 5258 16464 5264 16516
rect 5316 16504 5322 16516
rect 6825 16507 6883 16513
rect 6825 16504 6837 16507
rect 5316 16476 6837 16504
rect 5316 16464 5322 16476
rect 6825 16473 6837 16476
rect 6871 16473 6883 16507
rect 6825 16467 6883 16473
rect 7929 16507 7987 16513
rect 7929 16473 7941 16507
rect 7975 16504 7987 16507
rect 8478 16504 8484 16516
rect 7975 16476 8484 16504
rect 7975 16473 7987 16476
rect 7929 16467 7987 16473
rect 8478 16464 8484 16476
rect 8536 16464 8542 16516
rect 9227 16504 9255 16535
rect 9306 16532 9312 16584
rect 9364 16532 9370 16584
rect 9416 16581 9444 16612
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 13372 16640 13400 16671
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 13872 16680 14964 16708
rect 13872 16668 13878 16680
rect 14734 16640 14740 16652
rect 9861 16603 9919 16609
rect 11164 16612 12572 16640
rect 13372 16612 14740 16640
rect 9401 16575 9459 16581
rect 9401 16541 9413 16575
rect 9447 16541 9459 16575
rect 9401 16535 9459 16541
rect 9585 16575 9643 16581
rect 9585 16541 9597 16575
rect 9631 16572 9643 16575
rect 9674 16572 9680 16584
rect 9631 16544 9680 16572
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 11164 16581 11192 16612
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10192 16544 11161 16572
rect 10192 16532 10198 16544
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 11974 16572 11980 16584
rect 11149 16535 11207 16541
rect 11532 16544 11980 16572
rect 9227 16476 9674 16504
rect 5442 16436 5448 16448
rect 4908 16408 5448 16436
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6549 16439 6607 16445
rect 6549 16405 6561 16439
rect 6595 16436 6607 16439
rect 6638 16436 6644 16448
rect 6595 16408 6644 16436
rect 6595 16405 6607 16408
rect 6549 16399 6607 16405
rect 6638 16396 6644 16408
rect 6696 16396 6702 16448
rect 9025 16439 9083 16445
rect 9025 16405 9037 16439
rect 9071 16436 9083 16439
rect 9122 16436 9128 16448
rect 9071 16408 9128 16436
rect 9071 16405 9083 16408
rect 9025 16399 9083 16405
rect 9122 16396 9128 16408
rect 9180 16396 9186 16448
rect 9646 16436 9674 16476
rect 11054 16464 11060 16516
rect 11112 16504 11118 16516
rect 11532 16513 11560 16544
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12066 16532 12072 16584
rect 12124 16532 12130 16584
rect 12544 16581 12572 16612
rect 14734 16600 14740 16612
rect 14792 16600 14798 16652
rect 14936 16649 14964 16680
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15194 16640 15200 16652
rect 15151 16612 15200 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 15194 16600 15200 16612
rect 15252 16600 15258 16652
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 15804 16612 16497 16640
rect 15804 16600 15810 16612
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 12176 16544 12265 16572
rect 11517 16507 11575 16513
rect 11517 16504 11529 16507
rect 11112 16476 11529 16504
rect 11112 16464 11118 16476
rect 11517 16473 11529 16476
rect 11563 16473 11575 16507
rect 12176 16504 12204 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 12489 16575 12572 16581
rect 12489 16541 12501 16575
rect 12535 16544 12572 16575
rect 12535 16541 12547 16544
rect 12489 16535 12547 16541
rect 16022 16532 16028 16584
rect 16080 16572 16086 16584
rect 16393 16575 16451 16581
rect 16393 16572 16405 16575
rect 16080 16544 16405 16572
rect 16080 16532 16086 16544
rect 16393 16541 16405 16544
rect 16439 16541 16451 16575
rect 16393 16535 16451 16541
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 11517 16467 11575 16473
rect 11900 16476 12204 16504
rect 12345 16507 12403 16513
rect 10318 16436 10324 16448
rect 9646 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16436 10382 16448
rect 11900 16445 11928 16476
rect 12345 16473 12357 16507
rect 12391 16473 12403 16507
rect 12345 16467 12403 16473
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 10376 16408 11897 16436
rect 10376 16396 10382 16408
rect 11885 16405 11897 16408
rect 11931 16405 11943 16439
rect 11885 16399 11943 16405
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 12360 16436 12388 16467
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 14369 16507 14427 16513
rect 14369 16504 14381 16507
rect 13320 16476 14381 16504
rect 13320 16464 13326 16476
rect 14369 16473 14381 16476
rect 14415 16504 14427 16507
rect 15013 16507 15071 16513
rect 15013 16504 15025 16507
rect 14415 16476 15025 16504
rect 14415 16473 14427 16476
rect 14369 16467 14427 16473
rect 15013 16473 15025 16476
rect 15059 16473 15071 16507
rect 15013 16467 15071 16473
rect 12032 16408 12388 16436
rect 12032 16396 12038 16408
rect 12618 16396 12624 16448
rect 12676 16445 12682 16448
rect 12676 16399 12687 16445
rect 12676 16396 12682 16399
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 13538 16436 13544 16448
rect 13136 16408 13544 16436
rect 13136 16396 13142 16408
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 14550 16445 14556 16448
rect 14543 16439 14556 16445
rect 14543 16405 14555 16439
rect 14543 16399 14556 16405
rect 14550 16396 14556 16399
rect 14608 16396 14614 16448
rect 16850 16396 16856 16448
rect 16908 16396 16914 16448
rect 1104 16346 18860 16368
rect 1104 16294 3829 16346
rect 3881 16294 3893 16346
rect 3945 16294 3957 16346
rect 4009 16294 4021 16346
rect 4073 16294 4085 16346
rect 4137 16294 8268 16346
rect 8320 16294 8332 16346
rect 8384 16294 8396 16346
rect 8448 16294 8460 16346
rect 8512 16294 8524 16346
rect 8576 16294 12707 16346
rect 12759 16294 12771 16346
rect 12823 16294 12835 16346
rect 12887 16294 12899 16346
rect 12951 16294 12963 16346
rect 13015 16294 17146 16346
rect 17198 16294 17210 16346
rect 17262 16294 17274 16346
rect 17326 16294 17338 16346
rect 17390 16294 17402 16346
rect 17454 16294 18860 16346
rect 1104 16272 18860 16294
rect 5626 16232 5632 16244
rect 2976 16204 5632 16232
rect 2976 16108 3004 16204
rect 5626 16192 5632 16204
rect 5684 16192 5690 16244
rect 7101 16235 7159 16241
rect 7101 16201 7113 16235
rect 7147 16232 7159 16235
rect 10594 16232 10600 16244
rect 7147 16204 10600 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16201 12495 16235
rect 12437 16195 12495 16201
rect 4430 16164 4436 16176
rect 4370 16136 4436 16164
rect 4430 16124 4436 16136
rect 4488 16124 4494 16176
rect 9214 16164 9220 16176
rect 4632 16136 9220 16164
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 842 15988 848 16040
rect 900 16028 906 16040
rect 1581 16031 1639 16037
rect 1581 16028 1593 16031
rect 900 16000 1593 16028
rect 900 15988 906 16000
rect 1581 15997 1593 16000
rect 1627 15997 1639 16031
rect 1581 15991 1639 15997
rect 1872 15960 1900 16059
rect 2774 16056 2780 16108
rect 2832 16056 2838 16108
rect 2958 16056 2964 16108
rect 3016 16056 3022 16108
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 16028 2559 16031
rect 2590 16028 2596 16040
rect 2547 16000 2596 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 2590 15988 2596 16000
rect 2648 16028 2654 16040
rect 3234 16028 3240 16040
rect 2648 16000 3240 16028
rect 2648 15988 2654 16000
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 3329 16031 3387 16037
rect 3329 15997 3341 16031
rect 3375 16028 3387 16031
rect 4632 16028 4660 16136
rect 9214 16124 9220 16136
rect 9272 16124 9278 16176
rect 11790 16124 11796 16176
rect 11848 16164 11854 16176
rect 12069 16167 12127 16173
rect 12069 16164 12081 16167
rect 11848 16136 12081 16164
rect 11848 16124 11854 16136
rect 12069 16133 12081 16136
rect 12115 16133 12127 16167
rect 12452 16164 12480 16195
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 14093 16235 14151 16241
rect 14093 16232 14105 16235
rect 12584 16204 14105 16232
rect 12584 16192 12590 16204
rect 14093 16201 14105 16204
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 15378 16192 15384 16244
rect 15436 16192 15442 16244
rect 15562 16192 15568 16244
rect 15620 16192 15626 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 16666 16232 16672 16244
rect 16163 16204 16672 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 12452 16136 15332 16164
rect 12069 16127 12127 16133
rect 4706 16056 4712 16108
rect 4764 16096 4770 16108
rect 5902 16096 5908 16108
rect 4764 16068 5908 16096
rect 4764 16056 4770 16068
rect 5902 16056 5908 16068
rect 5960 16056 5966 16108
rect 6454 16056 6460 16108
rect 6512 16096 6518 16108
rect 8662 16105 8668 16108
rect 6733 16099 6791 16105
rect 6733 16096 6745 16099
rect 6512 16068 6745 16096
rect 6512 16056 6518 16068
rect 6733 16065 6745 16068
rect 6779 16065 6791 16099
rect 8660 16096 8668 16105
rect 8623 16068 8668 16096
rect 6733 16059 6791 16065
rect 8660 16059 8668 16068
rect 8662 16056 8668 16059
rect 8720 16056 8726 16108
rect 8754 16056 8760 16108
rect 8812 16056 8818 16108
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 9030 16096 9036 16108
rect 8956 16068 9036 16096
rect 3375 16000 4660 16028
rect 6549 16031 6607 16037
rect 3375 15997 3387 16000
rect 3329 15991 3387 15997
rect 6549 15997 6561 16031
rect 6595 15997 6607 16031
rect 6549 15991 6607 15997
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 6822 16028 6828 16040
rect 6687 16000 6828 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 6564 15960 6592 15991
rect 6822 15988 6828 16000
rect 6880 16028 6886 16040
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 6880 16000 7389 16028
rect 6880 15988 6886 16000
rect 7377 15997 7389 16000
rect 7423 15997 7435 16031
rect 7377 15991 7435 15997
rect 7929 16031 7987 16037
rect 7929 15997 7941 16031
rect 7975 16028 7987 16031
rect 8956 16028 8984 16068
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9122 16056 9128 16108
rect 9180 16056 9186 16108
rect 9646 16068 12664 16096
rect 7975 16000 8984 16028
rect 7975 15997 7987 16000
rect 7929 15991 7987 15997
rect 6914 15960 6920 15972
rect 1872 15932 3004 15960
rect 2976 15892 3004 15932
rect 4080 15932 5856 15960
rect 6564 15932 6920 15960
rect 4080 15892 4108 15932
rect 5828 15904 5856 15932
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7852 15932 8432 15960
rect 2976 15864 4108 15892
rect 5077 15895 5135 15901
rect 5077 15861 5089 15895
rect 5123 15892 5135 15895
rect 5166 15892 5172 15904
rect 5123 15864 5172 15892
rect 5123 15861 5135 15864
rect 5077 15855 5135 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5442 15852 5448 15904
rect 5500 15852 5506 15904
rect 5810 15852 5816 15904
rect 5868 15852 5874 15904
rect 7374 15852 7380 15904
rect 7432 15892 7438 15904
rect 7852 15892 7880 15932
rect 7432 15864 7880 15892
rect 7432 15852 7438 15864
rect 7926 15852 7932 15904
rect 7984 15892 7990 15904
rect 8202 15892 8208 15904
rect 7984 15864 8208 15892
rect 7984 15852 7990 15864
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 8404 15892 8432 15932
rect 8478 15920 8484 15972
rect 8536 15920 8542 15972
rect 8754 15920 8760 15972
rect 8812 15960 8818 15972
rect 9401 15963 9459 15969
rect 9401 15960 9413 15963
rect 8812 15932 9413 15960
rect 8812 15920 8818 15932
rect 9401 15929 9413 15932
rect 9447 15929 9459 15963
rect 9401 15923 9459 15929
rect 9646 15892 9674 16068
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 11664 16000 11805 16028
rect 11664 15988 11670 16000
rect 11793 15997 11805 16000
rect 11839 15997 11851 16031
rect 11793 15991 11851 15997
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 12636 16028 12664 16068
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 13538 16096 13544 16108
rect 13311 16068 13544 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 14274 16056 14280 16108
rect 14332 16056 14338 16108
rect 12986 16028 12992 16040
rect 12636 16000 12992 16028
rect 11977 15991 12035 15997
rect 11992 15960 12020 15991
rect 12986 15988 12992 16000
rect 13044 15988 13050 16040
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 15997 13139 16031
rect 15304 16028 15332 16136
rect 15396 16096 15424 16192
rect 15470 16124 15476 16176
rect 15528 16164 15534 16176
rect 16132 16164 16160 16195
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 15528 16136 16160 16164
rect 15528 16124 15534 16136
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15396 16068 15761 16096
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 17678 16028 17684 16040
rect 15304 16000 17684 16028
rect 13081 15991 13139 15997
rect 11256 15932 12020 15960
rect 11256 15904 11284 15932
rect 12526 15920 12532 15972
rect 12584 15920 12590 15972
rect 13096 15904 13124 15991
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 8404 15864 9674 15892
rect 9861 15895 9919 15901
rect 9861 15861 9873 15895
rect 9907 15892 9919 15895
rect 10318 15892 10324 15904
rect 9907 15864 10324 15892
rect 9907 15861 9919 15864
rect 9861 15855 9919 15861
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 11238 15852 11244 15904
rect 11296 15852 11302 15904
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 11882 15892 11888 15904
rect 11756 15864 11888 15892
rect 11756 15852 11762 15864
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 13078 15852 13084 15904
rect 13136 15892 13142 15904
rect 13633 15895 13691 15901
rect 13633 15892 13645 15895
rect 13136 15864 13645 15892
rect 13136 15852 13142 15864
rect 13633 15861 13645 15864
rect 13679 15861 13691 15895
rect 13633 15855 13691 15861
rect 1104 15802 18860 15824
rect 1104 15750 3169 15802
rect 3221 15750 3233 15802
rect 3285 15750 3297 15802
rect 3349 15750 3361 15802
rect 3413 15750 3425 15802
rect 3477 15750 7608 15802
rect 7660 15750 7672 15802
rect 7724 15750 7736 15802
rect 7788 15750 7800 15802
rect 7852 15750 7864 15802
rect 7916 15750 12047 15802
rect 12099 15750 12111 15802
rect 12163 15750 12175 15802
rect 12227 15750 12239 15802
rect 12291 15750 12303 15802
rect 12355 15750 16486 15802
rect 16538 15750 16550 15802
rect 16602 15750 16614 15802
rect 16666 15750 16678 15802
rect 16730 15750 16742 15802
rect 16794 15750 18860 15802
rect 1104 15728 18860 15750
rect 2225 15691 2283 15697
rect 2225 15657 2237 15691
rect 2271 15688 2283 15691
rect 2866 15688 2872 15700
rect 2271 15660 2872 15688
rect 2271 15657 2283 15660
rect 2225 15651 2283 15657
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 4341 15691 4399 15697
rect 4341 15688 4353 15691
rect 3568 15660 4353 15688
rect 3568 15648 3574 15660
rect 4341 15657 4353 15660
rect 4387 15657 4399 15691
rect 4341 15651 4399 15657
rect 5074 15648 5080 15700
rect 5132 15648 5138 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 6972 15660 7941 15688
rect 6972 15648 6978 15660
rect 7929 15657 7941 15660
rect 7975 15688 7987 15691
rect 7975 15660 12940 15688
rect 7975 15657 7987 15660
rect 7929 15651 7987 15657
rect 1581 15623 1639 15629
rect 1581 15589 1593 15623
rect 1627 15620 1639 15623
rect 10226 15620 10232 15632
rect 1627 15592 10232 15620
rect 1627 15589 1639 15592
rect 1581 15583 1639 15589
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 12912 15620 12940 15660
rect 12986 15648 12992 15700
rect 13044 15688 13050 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 13044 15660 17233 15688
rect 13044 15648 13050 15660
rect 17221 15657 17233 15660
rect 17267 15657 17279 15691
rect 17221 15651 17279 15657
rect 12912 15592 16988 15620
rect 1670 15512 1676 15564
rect 1728 15552 1734 15564
rect 2590 15552 2596 15564
rect 1728 15524 2596 15552
rect 1728 15512 1734 15524
rect 2590 15512 2596 15524
rect 2648 15552 2654 15564
rect 2869 15555 2927 15561
rect 2869 15552 2881 15555
rect 2648 15524 2881 15552
rect 2648 15512 2654 15524
rect 2869 15521 2881 15524
rect 2915 15521 2927 15555
rect 2869 15515 2927 15521
rect 6822 15512 6828 15564
rect 6880 15512 6886 15564
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15552 7251 15555
rect 7282 15552 7288 15564
rect 7239 15524 7288 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 7374 15512 7380 15564
rect 7432 15552 7438 15564
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 7432 15524 7481 15552
rect 7432 15512 7438 15524
rect 7469 15521 7481 15524
rect 7515 15521 7527 15555
rect 7469 15515 7527 15521
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 11238 15552 11244 15564
rect 8352 15524 11244 15552
rect 8352 15512 8358 15524
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11701 15555 11759 15561
rect 11701 15521 11713 15555
rect 11747 15552 11759 15555
rect 11882 15552 11888 15564
rect 11747 15524 11888 15552
rect 11747 15521 11759 15524
rect 11701 15515 11759 15521
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 11974 15512 11980 15564
rect 12032 15552 12038 15564
rect 16850 15552 16856 15564
rect 12032 15524 16856 15552
rect 12032 15512 12038 15524
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 1486 15444 1492 15496
rect 1544 15484 1550 15496
rect 3237 15487 3295 15493
rect 3237 15484 3249 15487
rect 1544 15456 3249 15484
rect 1544 15444 1550 15456
rect 3237 15453 3249 15456
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 3602 15444 3608 15496
rect 3660 15484 3666 15496
rect 4709 15487 4767 15493
rect 4709 15484 4721 15487
rect 3660 15456 4721 15484
rect 3660 15444 3666 15456
rect 4709 15453 4721 15456
rect 4755 15453 4767 15487
rect 4709 15447 4767 15453
rect 5810 15444 5816 15496
rect 5868 15484 5874 15496
rect 11330 15484 11336 15496
rect 5868 15456 11336 15484
rect 5868 15444 5874 15456
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 12066 15444 12072 15496
rect 12124 15444 12130 15496
rect 16960 15484 16988 15592
rect 17236 15552 17264 15651
rect 17236 15524 18184 15552
rect 17589 15487 17647 15493
rect 17589 15484 17601 15487
rect 16960 15456 17601 15484
rect 17589 15453 17601 15456
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 13084 15428 13136 15434
rect 2314 15376 2320 15428
rect 2372 15416 2378 15428
rect 2593 15419 2651 15425
rect 2593 15416 2605 15419
rect 2372 15388 2605 15416
rect 2372 15376 2378 15388
rect 2593 15385 2605 15388
rect 2639 15416 2651 15419
rect 3326 15416 3332 15428
rect 2639 15388 3332 15416
rect 2639 15385 2651 15388
rect 2593 15379 2651 15385
rect 3326 15376 3332 15388
rect 3384 15376 3390 15428
rect 4065 15419 4123 15425
rect 4065 15385 4077 15419
rect 4111 15416 4123 15419
rect 4246 15416 4252 15428
rect 4111 15388 4252 15416
rect 4111 15385 4123 15388
rect 4065 15379 4123 15385
rect 934 15308 940 15360
rect 992 15348 998 15360
rect 2406 15348 2412 15360
rect 992 15320 2412 15348
rect 992 15308 998 15320
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 3142 15308 3148 15360
rect 3200 15348 3206 15360
rect 4080 15348 4108 15379
rect 4246 15376 4252 15388
rect 4304 15416 4310 15428
rect 11238 15416 11244 15428
rect 4304 15388 11244 15416
rect 4304 15376 4310 15388
rect 11238 15376 11244 15388
rect 11296 15376 11302 15428
rect 13541 15419 13599 15425
rect 13541 15385 13553 15419
rect 13587 15416 13599 15419
rect 16390 15416 16396 15428
rect 13587 15388 16396 15416
rect 13587 15385 13599 15388
rect 13541 15379 13599 15385
rect 16390 15376 16396 15388
rect 16448 15376 16454 15428
rect 17604 15416 17632 15447
rect 17770 15444 17776 15496
rect 17828 15444 17834 15496
rect 17862 15444 17868 15496
rect 17920 15444 17926 15496
rect 18156 15493 18184 15524
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 18064 15416 18092 15447
rect 19242 15416 19248 15428
rect 17604 15388 19248 15416
rect 19242 15376 19248 15388
rect 19300 15376 19306 15428
rect 13084 15370 13136 15376
rect 3200 15320 4108 15348
rect 3200 15308 3206 15320
rect 4798 15308 4804 15360
rect 4856 15348 4862 15360
rect 8294 15348 8300 15360
rect 4856 15320 8300 15348
rect 4856 15308 4862 15320
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 8389 15351 8447 15357
rect 8389 15317 8401 15351
rect 8435 15348 8447 15351
rect 8662 15348 8668 15360
rect 8435 15320 8668 15348
rect 8435 15317 8447 15320
rect 8389 15311 8447 15317
rect 8662 15308 8668 15320
rect 8720 15348 8726 15360
rect 9950 15348 9956 15360
rect 8720 15320 9956 15348
rect 8720 15308 8726 15320
rect 9950 15308 9956 15320
rect 10008 15308 10014 15360
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11517 15351 11575 15357
rect 11517 15348 11529 15351
rect 10928 15320 11529 15348
rect 10928 15308 10934 15320
rect 11517 15317 11529 15320
rect 11563 15348 11575 15351
rect 11606 15348 11612 15360
rect 11563 15320 11612 15348
rect 11563 15317 11575 15320
rect 11517 15311 11575 15317
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 13909 15351 13967 15357
rect 13909 15317 13921 15351
rect 13955 15348 13967 15351
rect 14090 15348 14096 15360
rect 13955 15320 14096 15348
rect 13955 15317 13967 15320
rect 13909 15311 13967 15317
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 14642 15308 14648 15360
rect 14700 15308 14706 15360
rect 15010 15308 15016 15360
rect 15068 15308 15074 15360
rect 18322 15308 18328 15360
rect 18380 15308 18386 15360
rect 1104 15258 18860 15280
rect 1104 15206 3829 15258
rect 3881 15206 3893 15258
rect 3945 15206 3957 15258
rect 4009 15206 4021 15258
rect 4073 15206 4085 15258
rect 4137 15206 8268 15258
rect 8320 15206 8332 15258
rect 8384 15206 8396 15258
rect 8448 15206 8460 15258
rect 8512 15206 8524 15258
rect 8576 15206 12707 15258
rect 12759 15206 12771 15258
rect 12823 15206 12835 15258
rect 12887 15206 12899 15258
rect 12951 15206 12963 15258
rect 13015 15206 17146 15258
rect 17198 15206 17210 15258
rect 17262 15206 17274 15258
rect 17326 15206 17338 15258
rect 17390 15206 17402 15258
rect 17454 15206 18860 15258
rect 1104 15184 18860 15206
rect 1857 15147 1915 15153
rect 1857 15113 1869 15147
rect 1903 15144 1915 15147
rect 2314 15144 2320 15156
rect 1903 15116 2320 15144
rect 1903 15113 1915 15116
rect 1857 15107 1915 15113
rect 2314 15104 2320 15116
rect 2372 15104 2378 15156
rect 2958 15144 2964 15156
rect 2424 15116 2964 15144
rect 1486 14968 1492 15020
rect 1544 15008 1550 15020
rect 2424 15017 2452 15116
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 6454 15144 6460 15156
rect 3068 15116 6460 15144
rect 2774 15036 2780 15088
rect 2832 15076 2838 15088
rect 3068 15076 3096 15116
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 6822 15104 6828 15156
rect 6880 15144 6886 15156
rect 6880 15116 7420 15144
rect 6880 15104 6886 15116
rect 4430 15076 4436 15088
rect 2832 15048 3096 15076
rect 3910 15048 4436 15076
rect 2832 15036 2838 15048
rect 4430 15036 4436 15048
rect 4488 15076 4494 15088
rect 5718 15076 5724 15088
rect 4488 15048 5724 15076
rect 4488 15036 4494 15048
rect 5718 15036 5724 15048
rect 5776 15036 5782 15088
rect 5951 15079 6009 15085
rect 5951 15045 5963 15079
rect 5997 15076 6009 15079
rect 6546 15076 6552 15088
rect 5997 15048 6552 15076
rect 5997 15045 6009 15048
rect 5951 15039 6009 15045
rect 6546 15036 6552 15048
rect 6604 15036 6610 15088
rect 7282 15076 7288 15088
rect 6748 15048 7288 15076
rect 1765 15011 1823 15017
rect 1765 15008 1777 15011
rect 1544 14980 1777 15008
rect 1544 14968 1550 14980
rect 1765 14977 1777 14980
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 2409 15011 2467 15017
rect 2409 14977 2421 15011
rect 2455 14977 2467 15011
rect 4522 15008 4528 15020
rect 2409 14971 2467 14977
rect 3896 14980 4528 15008
rect 1670 14900 1676 14952
rect 1728 14900 1734 14952
rect 2682 14900 2688 14952
rect 2740 14900 2746 14952
rect 3326 14900 3332 14952
rect 3384 14940 3390 14952
rect 3896 14940 3924 14980
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 4982 14968 4988 15020
rect 5040 14968 5046 15020
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 14977 5227 15011
rect 5169 14971 5227 14977
rect 3384 14912 3924 14940
rect 3384 14900 3390 14912
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 4709 14943 4767 14949
rect 4709 14940 4721 14943
rect 4488 14912 4721 14940
rect 4488 14900 4494 14912
rect 4709 14909 4721 14912
rect 4755 14909 4767 14943
rect 4709 14903 4767 14909
rect 2038 14832 2044 14884
rect 2096 14872 2102 14884
rect 2406 14872 2412 14884
rect 2096 14844 2412 14872
rect 2096 14832 2102 14844
rect 2406 14832 2412 14844
rect 2464 14832 2470 14884
rect 4157 14875 4215 14881
rect 4157 14841 4169 14875
rect 4203 14872 4215 14875
rect 5074 14872 5080 14884
rect 4203 14844 5080 14872
rect 4203 14841 4215 14844
rect 4157 14835 4215 14841
rect 5074 14832 5080 14844
rect 5132 14832 5138 14884
rect 2225 14807 2283 14813
rect 2225 14773 2237 14807
rect 2271 14804 2283 14807
rect 4062 14804 4068 14816
rect 2271 14776 4068 14804
rect 2271 14773 2283 14776
rect 2225 14767 2283 14773
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4614 14764 4620 14816
rect 4672 14804 4678 14816
rect 5184 14804 5212 14971
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 5537 15011 5595 15017
rect 5537 15008 5549 15011
rect 5408 14980 5549 15008
rect 5408 14968 5414 14980
rect 5537 14977 5549 14980
rect 5583 15008 5595 15011
rect 6270 15008 6276 15020
rect 5583 14980 6276 15008
rect 5583 14977 5595 14980
rect 5537 14971 5595 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 6748 15017 6776 15048
rect 7282 15036 7288 15048
rect 7340 15036 7346 15088
rect 7392 15076 7420 15116
rect 8018 15104 8024 15156
rect 8076 15104 8082 15156
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 8386 15144 8392 15156
rect 8168 15116 8392 15144
rect 8168 15104 8174 15116
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 8588 15116 9168 15144
rect 8588 15076 8616 15116
rect 7392 15048 8616 15076
rect 9140 15076 9168 15116
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 9309 15147 9367 15153
rect 9309 15144 9321 15147
rect 9272 15116 9321 15144
rect 9272 15104 9278 15116
rect 9309 15113 9321 15116
rect 9355 15113 9367 15147
rect 9309 15107 9367 15113
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15344 15116 15945 15144
rect 15344 15104 15350 15116
rect 15933 15113 15945 15116
rect 15979 15144 15991 15147
rect 16206 15144 16212 15156
rect 15979 15116 16212 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 17770 15144 17776 15156
rect 17727 15116 17776 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 10410 15076 10416 15088
rect 9140 15048 10416 15076
rect 6640 15011 6698 15017
rect 6640 15008 6652 15011
rect 6380 14980 6652 15008
rect 5902 14900 5908 14952
rect 5960 14940 5966 14952
rect 6380 14940 6408 14980
rect 6640 14977 6652 14980
rect 6686 14977 6698 15011
rect 6640 14971 6698 14977
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 6914 15008 6920 15020
rect 6871 14980 6920 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 7392 15017 7420 15048
rect 10410 15036 10416 15048
rect 10468 15036 10474 15088
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 12253 15079 12311 15085
rect 12253 15076 12265 15079
rect 11480 15048 12265 15076
rect 11480 15036 11486 15048
rect 12253 15045 12265 15048
rect 12299 15045 12311 15079
rect 12253 15039 12311 15045
rect 12986 15036 12992 15088
rect 13044 15036 13050 15088
rect 14274 15036 14280 15088
rect 14332 15076 14338 15088
rect 16022 15076 16028 15088
rect 14332 15048 16028 15076
rect 14332 15036 14338 15048
rect 16022 15036 16028 15048
rect 16080 15036 16086 15088
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 15008 7067 15011
rect 7377 15011 7435 15017
rect 7055 14980 7328 15008
rect 7055 14977 7067 14980
rect 7009 14971 7067 14977
rect 7300 14952 7328 14980
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 5960 14912 6408 14940
rect 5960 14900 5966 14912
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 6512 14912 6961 14940
rect 6512 14900 6518 14912
rect 6365 14875 6423 14881
rect 6365 14841 6377 14875
rect 6411 14872 6423 14875
rect 6730 14872 6736 14884
rect 6411 14844 6736 14872
rect 6411 14841 6423 14844
rect 6365 14835 6423 14841
rect 6730 14832 6736 14844
rect 6788 14832 6794 14884
rect 4672 14776 5212 14804
rect 4672 14764 4678 14776
rect 5902 14764 5908 14816
rect 5960 14764 5966 14816
rect 6089 14807 6147 14813
rect 6089 14773 6101 14807
rect 6135 14804 6147 14807
rect 6454 14804 6460 14816
rect 6135 14776 6460 14804
rect 6135 14773 6147 14776
rect 6089 14767 6147 14773
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 6933 14804 6961 14912
rect 7282 14900 7288 14952
rect 7340 14900 7346 14952
rect 7466 14900 7472 14952
rect 7524 14900 7530 14952
rect 7760 14872 7788 14971
rect 8018 14968 8024 15020
rect 8076 14968 8082 15020
rect 8294 15016 8300 15020
rect 8266 15008 8300 15016
rect 8128 14980 8300 15008
rect 8128 14952 8156 14980
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 8570 14968 8576 15020
rect 8628 14998 8634 15020
rect 8665 15001 8723 15007
rect 8665 14998 8677 15001
rect 8628 14970 8677 14998
rect 8628 14968 8634 14970
rect 8665 14967 8677 14970
rect 8711 14967 8723 15001
rect 8846 14968 8852 15020
rect 8904 14968 8910 15020
rect 8938 14968 8944 15020
rect 8996 14968 9002 15020
rect 9214 14968 9220 15020
rect 9272 14968 9278 15020
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 15008 14427 15011
rect 15286 15008 15292 15020
rect 14415 14980 15292 15008
rect 14415 14977 14427 14980
rect 14369 14971 14427 14977
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 8665 14961 8723 14967
rect 8110 14900 8116 14952
rect 8168 14900 8174 14952
rect 8202 14900 8208 14952
rect 8260 14900 8266 14952
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 10042 14940 10048 14952
rect 9079 14912 10048 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 10042 14900 10048 14912
rect 10100 14900 10106 14952
rect 11882 14900 11888 14952
rect 11940 14940 11946 14952
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 11940 14912 11989 14940
rect 11940 14900 11946 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 11977 14903 12035 14909
rect 13648 14912 15577 14940
rect 10686 14872 10692 14884
rect 7760 14844 10692 14872
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 8478 14804 8484 14816
rect 6933 14776 8484 14804
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 8573 14807 8631 14813
rect 8573 14773 8585 14807
rect 8619 14804 8631 14807
rect 9214 14804 9220 14816
rect 8619 14776 9220 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 13648 14804 13676 14912
rect 15565 14909 15577 14912
rect 15611 14940 15623 14943
rect 16114 14940 16120 14952
rect 15611 14912 16120 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 14553 14875 14611 14881
rect 14553 14841 14565 14875
rect 14599 14872 14611 14875
rect 15010 14872 15016 14884
rect 14599 14844 15016 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 15010 14832 15016 14844
rect 15068 14832 15074 14884
rect 10560 14776 13676 14804
rect 10560 14764 10566 14776
rect 13722 14764 13728 14816
rect 13780 14764 13786 14816
rect 14001 14807 14059 14813
rect 14001 14773 14013 14807
rect 14047 14804 14059 14807
rect 14642 14804 14648 14816
rect 14047 14776 14648 14804
rect 14047 14773 14059 14776
rect 14001 14767 14059 14773
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 14918 14764 14924 14816
rect 14976 14764 14982 14816
rect 15286 14764 15292 14816
rect 15344 14804 15350 14816
rect 15930 14804 15936 14816
rect 15344 14776 15936 14804
rect 15344 14764 15350 14776
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 1104 14714 18860 14736
rect 1104 14662 3169 14714
rect 3221 14662 3233 14714
rect 3285 14662 3297 14714
rect 3349 14662 3361 14714
rect 3413 14662 3425 14714
rect 3477 14662 7608 14714
rect 7660 14662 7672 14714
rect 7724 14662 7736 14714
rect 7788 14662 7800 14714
rect 7852 14662 7864 14714
rect 7916 14662 12047 14714
rect 12099 14662 12111 14714
rect 12163 14662 12175 14714
rect 12227 14662 12239 14714
rect 12291 14662 12303 14714
rect 12355 14662 16486 14714
rect 16538 14662 16550 14714
rect 16602 14662 16614 14714
rect 16666 14662 16678 14714
rect 16730 14662 16742 14714
rect 16794 14662 18860 14714
rect 1104 14640 18860 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 3053 14603 3111 14609
rect 3053 14600 3065 14603
rect 1452 14572 3065 14600
rect 1452 14560 1458 14572
rect 3053 14569 3065 14572
rect 3099 14569 3111 14603
rect 3053 14563 3111 14569
rect 3513 14603 3571 14609
rect 3513 14569 3525 14603
rect 3559 14600 3571 14603
rect 4614 14600 4620 14612
rect 3559 14572 4620 14600
rect 3559 14569 3571 14572
rect 3513 14563 3571 14569
rect 1946 14492 1952 14544
rect 2004 14532 2010 14544
rect 3528 14532 3556 14563
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 5905 14603 5963 14609
rect 5905 14569 5917 14603
rect 5951 14600 5963 14603
rect 6178 14600 6184 14612
rect 5951 14572 6184 14600
rect 5951 14569 5963 14572
rect 5905 14563 5963 14569
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 7156 14572 7205 14600
rect 7156 14560 7162 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 7561 14603 7619 14609
rect 7561 14569 7573 14603
rect 7607 14600 7619 14603
rect 10962 14600 10968 14612
rect 7607 14572 10968 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11296 14572 14137 14600
rect 11296 14560 11302 14572
rect 2004 14504 3556 14532
rect 2004 14492 2010 14504
rect 7374 14492 7380 14544
rect 7432 14532 7438 14544
rect 7929 14535 7987 14541
rect 7929 14532 7941 14535
rect 7432 14504 7941 14532
rect 7432 14492 7438 14504
rect 7929 14501 7941 14504
rect 7975 14501 7987 14535
rect 8389 14535 8447 14541
rect 8389 14532 8401 14535
rect 7929 14495 7987 14501
rect 8266 14504 8401 14532
rect 1486 14424 1492 14476
rect 1544 14464 1550 14476
rect 2685 14467 2743 14473
rect 2685 14464 2697 14467
rect 1544 14436 2697 14464
rect 1544 14424 1550 14436
rect 2685 14433 2697 14436
rect 2731 14433 2743 14467
rect 2685 14427 2743 14433
rect 2958 14424 2964 14476
rect 3016 14464 3022 14476
rect 4157 14467 4215 14473
rect 4157 14464 4169 14467
rect 3016 14436 4169 14464
rect 3016 14424 3022 14436
rect 4157 14433 4169 14436
rect 4203 14433 4215 14467
rect 7392 14464 7420 14492
rect 4157 14427 4215 14433
rect 7208 14436 7420 14464
rect 1210 14356 1216 14408
rect 1268 14396 1274 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 1268 14368 1409 14396
rect 1268 14356 1274 14368
rect 1397 14365 1409 14368
rect 1443 14396 1455 14399
rect 2225 14399 2283 14405
rect 2225 14396 2237 14399
rect 1443 14368 2237 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2225 14365 2237 14368
rect 2271 14365 2283 14399
rect 5718 14396 5724 14408
rect 5566 14368 5724 14396
rect 2225 14359 2283 14365
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 6454 14356 6460 14408
rect 6512 14356 6518 14408
rect 7208 14405 7236 14436
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 7558 14396 7564 14408
rect 7423 14368 7564 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8266 14396 8294 14504
rect 8389 14501 8401 14504
rect 8435 14532 8447 14535
rect 8754 14532 8760 14544
rect 8435 14504 8760 14532
rect 8435 14501 8447 14504
rect 8389 14495 8447 14501
rect 8754 14492 8760 14504
rect 8812 14492 8818 14544
rect 8938 14492 8944 14544
rect 8996 14492 9002 14544
rect 13906 14532 13912 14544
rect 13464 14504 13912 14532
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 8956 14464 8984 14492
rect 8711 14436 8984 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 8168 14368 8294 14396
rect 8168 14356 8174 14368
rect 750 14288 756 14340
rect 808 14328 814 14340
rect 3970 14328 3976 14340
rect 808 14300 3976 14328
rect 808 14288 814 14300
rect 3970 14288 3976 14300
rect 4028 14288 4034 14340
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 4433 14331 4491 14337
rect 4433 14328 4445 14331
rect 4212 14300 4445 14328
rect 4212 14288 4218 14300
rect 4433 14297 4445 14300
rect 4479 14297 4491 14331
rect 6822 14328 6828 14340
rect 4433 14291 4491 14297
rect 5736 14300 6828 14328
rect 1578 14220 1584 14272
rect 1636 14220 1642 14272
rect 1670 14220 1676 14272
rect 1728 14260 1734 14272
rect 1857 14263 1915 14269
rect 1857 14260 1869 14263
rect 1728 14232 1869 14260
rect 1728 14220 1734 14232
rect 1857 14229 1869 14232
rect 1903 14229 1915 14263
rect 1857 14223 1915 14229
rect 4065 14263 4123 14269
rect 4065 14229 4077 14263
rect 4111 14260 4123 14263
rect 4338 14260 4344 14272
rect 4111 14232 4344 14260
rect 4111 14229 4123 14232
rect 4065 14223 4123 14229
rect 4338 14220 4344 14232
rect 4396 14260 4402 14272
rect 5736 14260 5764 14300
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 7576 14328 7604 14356
rect 8680 14328 8708 14427
rect 9306 14424 9312 14476
rect 9364 14424 9370 14476
rect 10134 14464 10140 14476
rect 9416 14436 10140 14464
rect 8938 14356 8944 14408
rect 8996 14356 9002 14408
rect 9416 14396 9444 14436
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 13464 14473 13492 14504
rect 13906 14492 13912 14504
rect 13964 14492 13970 14544
rect 14109 14532 14137 14572
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 14553 14603 14611 14609
rect 14553 14600 14565 14603
rect 14424 14572 14565 14600
rect 14424 14560 14430 14572
rect 14553 14569 14565 14572
rect 14599 14569 14611 14603
rect 14553 14563 14611 14569
rect 15013 14535 15071 14541
rect 15013 14532 15025 14535
rect 14109 14504 15025 14532
rect 15013 14501 15025 14504
rect 15059 14532 15071 14535
rect 15378 14532 15384 14544
rect 15059 14504 15384 14532
rect 15059 14501 15071 14504
rect 15013 14495 15071 14501
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 15657 14535 15715 14541
rect 15657 14501 15669 14535
rect 15703 14532 15715 14535
rect 19058 14532 19064 14544
rect 15703 14504 19064 14532
rect 15703 14501 15715 14504
rect 15657 14495 15715 14501
rect 19058 14492 19064 14504
rect 19116 14492 19122 14544
rect 13449 14467 13507 14473
rect 13449 14464 13461 14467
rect 11940 14436 13461 14464
rect 11940 14424 11946 14436
rect 13449 14433 13461 14436
rect 13495 14433 13507 14467
rect 13449 14427 13507 14433
rect 13740 14436 16068 14464
rect 9040 14368 9444 14396
rect 7576 14300 8708 14328
rect 4396 14232 5764 14260
rect 4396 14220 4402 14232
rect 6730 14220 6736 14272
rect 6788 14220 6794 14272
rect 6914 14220 6920 14272
rect 6972 14260 6978 14272
rect 9040 14260 9068 14368
rect 10778 14356 10784 14408
rect 10836 14356 10842 14408
rect 13740 14396 13768 14436
rect 13464 14368 13768 14396
rect 9582 14288 9588 14340
rect 9640 14328 9646 14340
rect 11517 14331 11575 14337
rect 9640 14300 9706 14328
rect 9640 14288 9646 14300
rect 11517 14297 11529 14331
rect 11563 14328 11575 14331
rect 13173 14331 13231 14337
rect 11563 14300 12006 14328
rect 11563 14297 11575 14300
rect 11517 14291 11575 14297
rect 6972 14232 9068 14260
rect 6972 14220 6978 14232
rect 9398 14220 9404 14272
rect 9456 14260 9462 14272
rect 9600 14260 9628 14288
rect 9456 14232 9628 14260
rect 9456 14220 9462 14232
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 11701 14263 11759 14269
rect 11701 14260 11713 14263
rect 10192 14232 11713 14260
rect 10192 14220 10198 14232
rect 11701 14229 11713 14232
rect 11747 14229 11759 14263
rect 11900 14260 11928 14300
rect 13173 14297 13185 14331
rect 13219 14328 13231 14331
rect 13464 14328 13492 14368
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13872 14368 14105 14396
rect 13872 14356 13878 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14366 14356 14372 14408
rect 14424 14356 14430 14408
rect 15562 14356 15568 14408
rect 15620 14356 15626 14408
rect 16040 14396 16068 14436
rect 16114 14424 16120 14476
rect 16172 14424 16178 14476
rect 16206 14424 16212 14476
rect 16264 14424 16270 14476
rect 19150 14396 19156 14408
rect 16040 14368 19156 14396
rect 19150 14356 19156 14368
rect 19208 14356 19214 14408
rect 13219 14300 13492 14328
rect 13648 14300 14228 14328
rect 13219 14297 13231 14300
rect 13173 14291 13231 14297
rect 12526 14260 12532 14272
rect 11900 14232 12532 14260
rect 11701 14223 11759 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 13648 14260 13676 14300
rect 13412 14232 13676 14260
rect 13412 14220 13418 14232
rect 13814 14220 13820 14272
rect 13872 14220 13878 14272
rect 14200 14269 14228 14300
rect 14274 14288 14280 14340
rect 14332 14328 14338 14340
rect 16298 14328 16304 14340
rect 14332 14300 16304 14328
rect 14332 14288 14338 14300
rect 16298 14288 16304 14300
rect 16356 14288 16362 14340
rect 14185 14263 14243 14269
rect 14185 14229 14197 14263
rect 14231 14229 14243 14263
rect 14185 14223 14243 14229
rect 15381 14263 15439 14269
rect 15381 14229 15393 14263
rect 15427 14260 15439 14263
rect 15654 14260 15660 14272
rect 15427 14232 15660 14260
rect 15427 14229 15439 14232
rect 15381 14223 15439 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 16025 14263 16083 14269
rect 16025 14260 16037 14263
rect 15896 14232 16037 14260
rect 15896 14220 15902 14232
rect 16025 14229 16037 14232
rect 16071 14229 16083 14263
rect 16025 14223 16083 14229
rect 1104 14170 18860 14192
rect 1104 14118 3829 14170
rect 3881 14118 3893 14170
rect 3945 14118 3957 14170
rect 4009 14118 4021 14170
rect 4073 14118 4085 14170
rect 4137 14118 8268 14170
rect 8320 14118 8332 14170
rect 8384 14118 8396 14170
rect 8448 14118 8460 14170
rect 8512 14118 8524 14170
rect 8576 14118 12707 14170
rect 12759 14118 12771 14170
rect 12823 14118 12835 14170
rect 12887 14118 12899 14170
rect 12951 14118 12963 14170
rect 13015 14118 17146 14170
rect 17198 14118 17210 14170
rect 17262 14118 17274 14170
rect 17326 14118 17338 14170
rect 17390 14118 17402 14170
rect 17454 14118 18860 14170
rect 1104 14096 18860 14118
rect 1578 14016 1584 14068
rect 1636 14016 1642 14068
rect 5350 14056 5356 14068
rect 4080 14028 5356 14056
rect 3694 13988 3700 14000
rect 3528 13960 3700 13988
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 2777 13923 2835 13929
rect 2777 13920 2789 13923
rect 1452 13892 2789 13920
rect 1452 13880 1458 13892
rect 2777 13889 2789 13892
rect 2823 13889 2835 13923
rect 2777 13883 2835 13889
rect 3050 13880 3056 13932
rect 3108 13920 3114 13932
rect 3528 13929 3556 13960
rect 3694 13948 3700 13960
rect 3752 13948 3758 14000
rect 4080 13929 4108 14028
rect 5350 14016 5356 14028
rect 5408 14056 5414 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 5408 14028 5733 14056
rect 5408 14016 5414 14028
rect 5721 14025 5733 14028
rect 5767 14056 5779 14059
rect 8018 14056 8024 14068
rect 5767 14028 8024 14056
rect 5767 14025 5779 14028
rect 5721 14019 5779 14025
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 12618 14056 12624 14068
rect 11388 14028 12624 14056
rect 11388 14016 11394 14028
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 13538 14056 13544 14068
rect 13044 14028 13544 14056
rect 13044 14016 13050 14028
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 13998 14056 14004 14068
rect 13648 14028 14004 14056
rect 4433 13991 4491 13997
rect 4433 13957 4445 13991
rect 4479 13988 4491 13991
rect 4479 13960 5120 13988
rect 4479 13957 4491 13960
rect 4433 13951 4491 13957
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 3108 13892 3249 13920
rect 3108 13880 3114 13892
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 4065 13923 4123 13929
rect 4065 13889 4077 13923
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 4338 13880 4344 13932
rect 4396 13880 4402 13932
rect 4571 13923 4629 13929
rect 4571 13889 4583 13923
rect 4617 13920 4629 13923
rect 5092 13920 5120 13960
rect 6086 13948 6092 14000
rect 6144 13988 6150 14000
rect 6914 13988 6920 14000
rect 6144 13960 6920 13988
rect 6144 13948 6150 13960
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 7745 13991 7803 13997
rect 7745 13988 7757 13991
rect 7156 13960 7757 13988
rect 7156 13948 7162 13960
rect 7745 13957 7757 13960
rect 7791 13957 7803 13991
rect 7745 13951 7803 13957
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 9364 13960 9812 13988
rect 9364 13948 9370 13960
rect 4617 13892 5028 13920
rect 5092 13892 5212 13920
rect 4617 13889 4629 13892
rect 4571 13883 4629 13889
rect 2038 13812 2044 13864
rect 2096 13812 2102 13864
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 2924 13824 3341 13852
rect 2924 13812 2930 13824
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 3329 13815 3387 13821
rect 3970 13812 3976 13864
rect 4028 13812 4034 13864
rect 4586 13852 4614 13883
rect 4890 13852 4896 13864
rect 4172 13824 4614 13852
rect 4724 13824 4896 13852
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 2409 13719 2467 13725
rect 2409 13716 2421 13719
rect 2004 13688 2421 13716
rect 2004 13676 2010 13688
rect 2409 13685 2421 13688
rect 2455 13685 2467 13719
rect 2409 13679 2467 13685
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 4172 13716 4200 13824
rect 4724 13725 4752 13824
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5000 13784 5028 13892
rect 5184 13852 5212 13892
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 9398 13920 9404 13932
rect 7524 13892 9404 13920
rect 7524 13880 7530 13892
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13889 9551 13923
rect 9784 13923 9812 13960
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 13648 13988 13676 14028
rect 13998 14016 14004 14028
rect 14056 14056 14062 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 14056 14028 14473 14056
rect 14056 14016 14062 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 16264 14028 16865 14056
rect 16264 14016 16270 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 10008 13960 13676 13988
rect 10008 13948 10014 13960
rect 14090 13948 14096 14000
rect 14148 13948 14154 14000
rect 14550 13948 14556 14000
rect 14608 13988 14614 14000
rect 14608 13960 15410 13988
rect 14608 13948 14614 13960
rect 9862 13926 9920 13932
rect 9862 13923 9874 13926
rect 9784 13895 9874 13923
rect 9493 13883 9551 13889
rect 9862 13892 9874 13895
rect 9908 13892 9920 13926
rect 9862 13886 9920 13892
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13918 10103 13923
rect 10226 13920 10232 13932
rect 10152 13918 10232 13920
rect 10091 13892 10232 13918
rect 10091 13890 10180 13892
rect 10091 13889 10103 13890
rect 10045 13883 10103 13889
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 5184 13824 5365 13852
rect 5353 13821 5365 13824
rect 5399 13852 5411 13855
rect 7006 13852 7012 13864
rect 5399 13824 7012 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 9309 13855 9367 13861
rect 9309 13852 9321 13855
rect 8720 13824 9321 13852
rect 8720 13812 8726 13824
rect 9309 13821 9321 13824
rect 9355 13821 9367 13855
rect 9309 13815 9367 13821
rect 6086 13784 6092 13796
rect 5000 13756 6092 13784
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 7098 13744 7104 13796
rect 7156 13784 7162 13796
rect 9214 13784 9220 13796
rect 7156 13756 9220 13784
rect 7156 13744 7162 13756
rect 9214 13744 9220 13756
rect 9272 13784 9278 13796
rect 9508 13784 9536 13883
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 10410 13880 10416 13932
rect 10468 13920 10474 13932
rect 10468 13892 12480 13920
rect 10468 13880 10474 13892
rect 9674 13812 9680 13864
rect 9732 13812 9738 13864
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 12452 13852 12480 13892
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 12986 13920 12992 13932
rect 12584 13892 12992 13920
rect 12584 13880 12590 13892
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 13630 13852 13636 13864
rect 9824 13824 10456 13852
rect 12452 13824 13636 13852
rect 9824 13812 9830 13824
rect 10428 13793 10456 13824
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14458 13852 14464 13864
rect 13964 13824 14464 13852
rect 13964 13812 13970 13824
rect 14458 13812 14464 13824
rect 14516 13852 14522 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14516 13824 14657 13852
rect 14516 13812 14522 13824
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 14918 13812 14924 13864
rect 14976 13812 14982 13864
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 16298 13852 16304 13864
rect 15068 13824 16304 13852
rect 15068 13812 15074 13824
rect 16298 13812 16304 13824
rect 16356 13852 16362 13864
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 16356 13824 16405 13852
rect 16356 13812 16362 13824
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 10413 13787 10471 13793
rect 9272 13756 9904 13784
rect 9272 13744 9278 13756
rect 2648 13688 4200 13716
rect 4709 13719 4767 13725
rect 2648 13676 2654 13688
rect 4709 13685 4721 13719
rect 4755 13685 4767 13719
rect 4709 13679 4767 13685
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 7009 13719 7067 13725
rect 7009 13716 7021 13719
rect 5224 13688 7021 13716
rect 5224 13676 5230 13688
rect 7009 13685 7021 13688
rect 7055 13716 7067 13719
rect 7466 13716 7472 13728
rect 7055 13688 7472 13716
rect 7055 13685 7067 13688
rect 7009 13679 7067 13685
rect 7466 13676 7472 13688
rect 7524 13676 7530 13728
rect 8849 13719 8907 13725
rect 8849 13685 8861 13719
rect 8895 13716 8907 13719
rect 9306 13716 9312 13728
rect 8895 13688 9312 13716
rect 8895 13685 8907 13688
rect 8849 13679 8907 13685
rect 9306 13676 9312 13688
rect 9364 13676 9370 13728
rect 9876 13716 9904 13756
rect 10413 13753 10425 13787
rect 10459 13784 10471 13787
rect 10778 13784 10784 13796
rect 10459 13756 10784 13784
rect 10459 13753 10471 13756
rect 10413 13747 10471 13753
rect 10778 13744 10784 13756
rect 10836 13784 10842 13796
rect 14274 13784 14280 13796
rect 10836 13756 14280 13784
rect 10836 13744 10842 13756
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 11793 13719 11851 13725
rect 11793 13716 11805 13719
rect 9876 13688 11805 13716
rect 11793 13685 11805 13688
rect 11839 13716 11851 13719
rect 11882 13716 11888 13728
rect 11839 13688 11888 13716
rect 11839 13685 11851 13688
rect 11793 13679 11851 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13722 13716 13728 13728
rect 13136 13688 13728 13716
rect 13136 13676 13142 13688
rect 13722 13676 13728 13688
rect 13780 13676 13786 13728
rect 1104 13626 18860 13648
rect 1104 13574 3169 13626
rect 3221 13574 3233 13626
rect 3285 13574 3297 13626
rect 3349 13574 3361 13626
rect 3413 13574 3425 13626
rect 3477 13574 7608 13626
rect 7660 13574 7672 13626
rect 7724 13574 7736 13626
rect 7788 13574 7800 13626
rect 7852 13574 7864 13626
rect 7916 13574 12047 13626
rect 12099 13574 12111 13626
rect 12163 13574 12175 13626
rect 12227 13574 12239 13626
rect 12291 13574 12303 13626
rect 12355 13574 16486 13626
rect 16538 13574 16550 13626
rect 16602 13574 16614 13626
rect 16666 13574 16678 13626
rect 16730 13574 16742 13626
rect 16794 13574 18860 13626
rect 1104 13552 18860 13574
rect 2133 13515 2191 13521
rect 2133 13481 2145 13515
rect 2179 13512 2191 13515
rect 2498 13512 2504 13524
rect 2179 13484 2504 13512
rect 2179 13481 2191 13484
rect 2133 13475 2191 13481
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 4430 13512 4436 13524
rect 4120 13484 4436 13512
rect 4120 13472 4126 13484
rect 4430 13472 4436 13484
rect 4488 13472 4494 13524
rect 9950 13512 9956 13524
rect 5000 13484 9956 13512
rect 5000 13444 5028 13484
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 13262 13512 13268 13524
rect 10468 13484 13268 13512
rect 10468 13472 10474 13484
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 13630 13472 13636 13524
rect 13688 13472 13694 13524
rect 13722 13472 13728 13524
rect 13780 13512 13786 13524
rect 13906 13512 13912 13524
rect 13780 13484 13912 13512
rect 13780 13472 13786 13484
rect 13906 13472 13912 13484
rect 13964 13512 13970 13524
rect 14277 13515 14335 13521
rect 14277 13512 14289 13515
rect 13964 13484 14289 13512
rect 13964 13472 13970 13484
rect 14277 13481 14289 13484
rect 14323 13481 14335 13515
rect 15194 13512 15200 13524
rect 14277 13475 14335 13481
rect 14383 13484 15200 13512
rect 4264 13416 5028 13444
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13376 2927 13379
rect 4154 13376 4160 13388
rect 2915 13348 4160 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 4154 13336 4160 13348
rect 4212 13336 4218 13388
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1670 13308 1676 13320
rect 1452 13280 1676 13308
rect 1452 13268 1458 13280
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 1854 13268 1860 13320
rect 1912 13268 1918 13320
rect 1946 13268 1952 13320
rect 2004 13268 2010 13320
rect 3142 13268 3148 13320
rect 3200 13308 3206 13320
rect 3694 13308 3700 13320
rect 3200 13280 3700 13308
rect 3200 13268 3206 13280
rect 3694 13268 3700 13280
rect 3752 13268 3758 13320
rect 4264 13317 4292 13416
rect 7466 13404 7472 13456
rect 7524 13444 7530 13456
rect 7837 13447 7895 13453
rect 7837 13444 7849 13447
rect 7524 13416 7849 13444
rect 7524 13404 7530 13416
rect 7837 13413 7849 13416
rect 7883 13413 7895 13447
rect 7837 13407 7895 13413
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 8168 13416 8294 13444
rect 8168 13404 8174 13416
rect 4522 13336 4528 13388
rect 4580 13336 4586 13388
rect 6270 13336 6276 13388
rect 6328 13336 6334 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 8018 13376 8024 13388
rect 7708 13348 8024 13376
rect 7708 13336 7714 13348
rect 8018 13336 8024 13348
rect 8076 13336 8082 13388
rect 8266 13376 8294 13416
rect 11882 13404 11888 13456
rect 11940 13444 11946 13456
rect 12250 13444 12256 13456
rect 11940 13416 12256 13444
rect 11940 13404 11946 13416
rect 12250 13404 12256 13416
rect 12308 13444 12314 13456
rect 12308 13416 12480 13444
rect 12308 13404 12314 13416
rect 11609 13379 11667 13385
rect 11609 13376 11621 13379
rect 8266 13348 11621 13376
rect 11609 13345 11621 13348
rect 11655 13376 11667 13379
rect 12452 13376 12480 13416
rect 12894 13404 12900 13456
rect 12952 13444 12958 13456
rect 13357 13447 13415 13453
rect 13357 13444 13369 13447
rect 12952 13416 13369 13444
rect 12952 13404 12958 13416
rect 13357 13413 13369 13416
rect 13403 13444 13415 13447
rect 14383 13444 14411 13484
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 16022 13512 16028 13524
rect 15436 13484 16028 13512
rect 15436 13472 15442 13484
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 16209 13447 16267 13453
rect 13403 13416 14411 13444
rect 14476 13416 15700 13444
rect 13403 13413 13415 13416
rect 13357 13407 13415 13413
rect 14476 13376 14504 13416
rect 11655 13348 12388 13376
rect 12452 13348 14504 13376
rect 11655 13345 11667 13348
rect 11609 13339 11667 13345
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 9674 13308 9680 13320
rect 6788 13280 9680 13308
rect 6788 13268 6794 13280
rect 9674 13268 9680 13280
rect 9732 13308 9738 13320
rect 10870 13308 10876 13320
rect 9732 13280 10876 13308
rect 9732 13268 9738 13280
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 10962 13268 10968 13320
rect 11020 13308 11026 13320
rect 11881 13317 11909 13348
rect 11701 13311 11759 13317
rect 11701 13308 11713 13311
rect 11020 13280 11713 13308
rect 11020 13268 11026 13280
rect 11701 13277 11713 13280
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 11866 13311 11924 13317
rect 11866 13277 11878 13311
rect 11912 13308 11924 13311
rect 11977 13311 12035 13317
rect 11912 13280 11946 13308
rect 11912 13277 11924 13280
rect 11866 13271 11924 13277
rect 11977 13277 11989 13311
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 1596 13212 2774 13240
rect 1596 13181 1624 13212
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 1762 13172 1768 13184
rect 1719 13144 1768 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 2314 13172 2320 13184
rect 1912 13144 2320 13172
rect 1912 13132 1918 13144
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 2406 13132 2412 13184
rect 2464 13172 2470 13184
rect 2501 13175 2559 13181
rect 2501 13172 2513 13175
rect 2464 13144 2513 13172
rect 2464 13132 2470 13144
rect 2501 13141 2513 13144
rect 2547 13172 2559 13175
rect 2590 13172 2596 13184
rect 2547 13144 2596 13172
rect 2547 13141 2559 13144
rect 2501 13135 2559 13141
rect 2590 13132 2596 13144
rect 2648 13132 2654 13184
rect 2746 13172 2774 13212
rect 3602 13200 3608 13252
rect 3660 13200 3666 13252
rect 3973 13243 4031 13249
rect 3973 13209 3985 13243
rect 4019 13240 4031 13243
rect 4706 13240 4712 13252
rect 4019 13212 4712 13240
rect 4019 13209 4031 13212
rect 3973 13203 4031 13209
rect 4706 13200 4712 13212
rect 4764 13200 4770 13252
rect 5718 13240 5724 13252
rect 5566 13212 5724 13240
rect 5718 13200 5724 13212
rect 5776 13200 5782 13252
rect 5994 13200 6000 13252
rect 6052 13200 6058 13252
rect 6086 13200 6092 13252
rect 6144 13240 6150 13252
rect 10134 13240 10140 13252
rect 6144 13212 10140 13240
rect 6144 13200 6150 13212
rect 10134 13200 10140 13212
rect 10192 13200 10198 13252
rect 11238 13200 11244 13252
rect 11296 13200 11302 13252
rect 11330 13200 11336 13252
rect 11388 13240 11394 13252
rect 11992 13240 12020 13271
rect 12066 13268 12072 13320
rect 12124 13268 12130 13320
rect 12250 13268 12256 13320
rect 12308 13268 12314 13320
rect 12360 13308 12388 13348
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 15010 13376 15016 13388
rect 14792 13348 15016 13376
rect 14792 13336 14798 13348
rect 15010 13336 15016 13348
rect 15068 13336 15074 13388
rect 15378 13336 15384 13388
rect 15436 13336 15442 13388
rect 12360 13280 13124 13308
rect 12713 13243 12771 13249
rect 12713 13240 12725 13243
rect 11388 13212 12725 13240
rect 11388 13200 11394 13212
rect 12713 13209 12725 13212
rect 12759 13209 12771 13243
rect 13096 13240 13124 13280
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 15105 13311 15163 13317
rect 15105 13308 15117 13311
rect 13504 13280 15117 13308
rect 13504 13268 13510 13280
rect 15105 13277 15117 13280
rect 15151 13277 15163 13311
rect 15286 13308 15292 13320
rect 15247 13280 15292 13308
rect 15105 13271 15163 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15672 13317 15700 13416
rect 16209 13413 16221 13447
rect 16255 13444 16267 13447
rect 18598 13444 18604 13456
rect 16255 13416 18604 13444
rect 16255 13413 16267 13416
rect 16209 13407 16267 13413
rect 18598 13404 18604 13416
rect 18656 13404 18662 13456
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 15804 13348 17049 13376
rect 15804 13336 15810 13348
rect 17037 13345 17049 13348
rect 17083 13345 17095 13379
rect 17037 13339 17095 13345
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 16393 13311 16451 13317
rect 15703 13280 15884 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 13538 13240 13544 13252
rect 13096 13212 13544 13240
rect 12713 13203 12771 13209
rect 13538 13200 13544 13212
rect 13596 13200 13602 13252
rect 14090 13200 14096 13252
rect 14148 13240 14154 13252
rect 14274 13240 14280 13252
rect 14148 13212 14280 13240
rect 14148 13200 14154 13212
rect 14274 13200 14280 13212
rect 14332 13240 14338 13252
rect 15488 13240 15516 13271
rect 14332 13212 15516 13240
rect 14332 13200 14338 13212
rect 5074 13172 5080 13184
rect 2746 13144 5080 13172
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5626 13132 5632 13184
rect 5684 13172 5690 13184
rect 6730 13172 6736 13184
rect 5684 13144 6736 13172
rect 5684 13132 5690 13144
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 9122 13132 9128 13184
rect 9180 13132 9186 13184
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9456 13144 9505 13172
rect 9456 13132 9462 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 11882 13172 11888 13184
rect 9824 13144 11888 13172
rect 9824 13132 9830 13144
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 12345 13175 12403 13181
rect 12345 13141 12357 13175
rect 12391 13172 12403 13175
rect 13446 13172 13452 13184
rect 12391 13144 13452 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 13446 13132 13452 13144
rect 13504 13132 13510 13184
rect 14918 13132 14924 13184
rect 14976 13172 14982 13184
rect 15749 13175 15807 13181
rect 15749 13172 15761 13175
rect 14976 13144 15761 13172
rect 14976 13132 14982 13144
rect 15749 13141 15761 13144
rect 15795 13141 15807 13175
rect 15856 13172 15884 13280
rect 16393 13277 16405 13311
rect 16439 13308 16451 13311
rect 16482 13308 16488 13320
rect 16439 13280 16488 13308
rect 16439 13277 16451 13280
rect 16393 13271 16451 13277
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 16666 13200 16672 13252
rect 16724 13200 16730 13252
rect 17497 13175 17555 13181
rect 17497 13172 17509 13175
rect 15856 13144 17509 13172
rect 15749 13135 15807 13141
rect 17497 13141 17509 13144
rect 17543 13172 17555 13175
rect 17586 13172 17592 13184
rect 17543 13144 17592 13172
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 1104 13082 18860 13104
rect 1104 13030 3829 13082
rect 3881 13030 3893 13082
rect 3945 13030 3957 13082
rect 4009 13030 4021 13082
rect 4073 13030 4085 13082
rect 4137 13030 8268 13082
rect 8320 13030 8332 13082
rect 8384 13030 8396 13082
rect 8448 13030 8460 13082
rect 8512 13030 8524 13082
rect 8576 13030 12707 13082
rect 12759 13030 12771 13082
rect 12823 13030 12835 13082
rect 12887 13030 12899 13082
rect 12951 13030 12963 13082
rect 13015 13030 17146 13082
rect 17198 13030 17210 13082
rect 17262 13030 17274 13082
rect 17326 13030 17338 13082
rect 17390 13030 17402 13082
rect 17454 13030 18860 13082
rect 1104 13008 18860 13030
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 3418 12968 3424 12980
rect 3016 12940 3424 12968
rect 3016 12928 3022 12940
rect 3418 12928 3424 12940
rect 3476 12928 3482 12980
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 9122 12968 9128 12980
rect 3844 12940 9128 12968
rect 3844 12928 3850 12940
rect 5261 12903 5319 12909
rect 2898 12886 3556 12900
rect 2884 12872 3556 12886
rect 4830 12872 4936 12900
rect 1489 12835 1547 12841
rect 1489 12801 1501 12835
rect 1535 12832 1547 12835
rect 1535 12804 1992 12832
rect 1535 12801 1547 12804
rect 1489 12795 1547 12801
rect 1854 12724 1860 12776
rect 1912 12724 1918 12776
rect 1964 12764 1992 12804
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 2884 12832 2912 12872
rect 3418 12832 3424 12844
rect 2740 12804 2912 12832
rect 2976 12804 3424 12832
rect 2740 12792 2746 12804
rect 2976 12764 3004 12804
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 3528 12832 3556 12872
rect 3528 12804 3924 12832
rect 3789 12767 3847 12773
rect 3789 12764 3801 12767
rect 1964 12736 3004 12764
rect 3068 12736 3801 12764
rect 1026 12588 1032 12640
rect 1084 12628 1090 12640
rect 3068 12628 3096 12736
rect 3789 12733 3801 12736
rect 3835 12733 3847 12767
rect 3896 12764 3924 12804
rect 4908 12764 4936 12872
rect 5261 12869 5273 12903
rect 5307 12900 5319 12903
rect 7650 12900 7656 12912
rect 5307 12872 7656 12900
rect 5307 12869 5319 12872
rect 5261 12863 5319 12869
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 8496 12909 8524 12940
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 9263 12940 9965 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 9953 12937 9965 12940
rect 9999 12968 10011 12971
rect 10410 12968 10416 12980
rect 9999 12940 10416 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 7929 12903 7987 12909
rect 7929 12869 7941 12903
rect 7975 12900 7987 12903
rect 8389 12903 8447 12909
rect 8389 12900 8401 12903
rect 7975 12872 8401 12900
rect 7975 12869 7987 12872
rect 7929 12863 7987 12869
rect 8389 12869 8401 12872
rect 8435 12869 8447 12903
rect 8389 12863 8447 12869
rect 8481 12903 8539 12909
rect 8481 12869 8493 12903
rect 8527 12869 8539 12903
rect 8846 12900 8852 12912
rect 8481 12863 8539 12869
rect 8588 12872 8852 12900
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5224 12804 5641 12832
rect 5224 12792 5230 12804
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 6178 12832 6184 12844
rect 5767 12804 6184 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 3896 12736 4936 12764
rect 3789 12727 3847 12733
rect 1084 12600 3096 12628
rect 3237 12631 3295 12637
rect 1084 12588 1090 12600
rect 3237 12597 3249 12631
rect 3283 12628 3295 12631
rect 3694 12628 3700 12640
rect 3283 12600 3700 12628
rect 3283 12597 3295 12600
rect 3237 12591 3295 12597
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4614 12628 4620 12640
rect 4212 12600 4620 12628
rect 4212 12588 4218 12600
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 4908 12628 4936 12736
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 5644 12764 5672 12795
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 7944 12832 7972 12863
rect 8294 12841 8300 12844
rect 8292 12832 8300 12841
rect 6512 12804 7972 12832
rect 8255 12804 8300 12832
rect 6512 12792 6518 12804
rect 8292 12795 8300 12804
rect 8294 12792 8300 12795
rect 8352 12792 8358 12844
rect 8404 12832 8432 12863
rect 8588 12832 8616 12872
rect 8846 12860 8852 12872
rect 8904 12860 8910 12912
rect 8938 12860 8944 12912
rect 8996 12900 9002 12912
rect 9232 12900 9260 12931
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 12158 12968 12164 12980
rect 11204 12940 12164 12968
rect 11204 12928 11210 12940
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12250 12928 12256 12980
rect 12308 12968 12314 12980
rect 12802 12968 12808 12980
rect 12308 12940 12808 12968
rect 12308 12928 12314 12940
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 13722 12968 13728 12980
rect 13556 12940 13728 12968
rect 8996 12872 9260 12900
rect 10045 12903 10103 12909
rect 8996 12860 9002 12872
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 10870 12900 10876 12912
rect 10091 12872 10876 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 8404 12804 8616 12832
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9674 12832 9680 12844
rect 9631 12804 9680 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 5644 12736 6929 12764
rect 5537 12727 5595 12733
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 5552 12696 5580 12727
rect 6932 12696 6960 12727
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 8680 12764 8708 12795
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 10060 12832 10088 12863
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 13556 12900 13584 12940
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12968 13967 12971
rect 14182 12968 14188 12980
rect 13955 12940 14188 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 15470 12968 15476 12980
rect 14384 12940 15476 12968
rect 13202 12872 13584 12900
rect 13630 12860 13636 12912
rect 13688 12900 13694 12912
rect 14384 12909 14412 12940
rect 15470 12928 15476 12940
rect 15528 12968 15534 12980
rect 15838 12968 15844 12980
rect 15528 12940 15844 12968
rect 15528 12928 15534 12940
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 15933 12971 15991 12977
rect 15933 12937 15945 12971
rect 15979 12968 15991 12971
rect 16390 12968 16396 12980
rect 15979 12940 16396 12968
rect 15979 12937 15991 12940
rect 15933 12931 15991 12937
rect 16390 12928 16396 12940
rect 16448 12968 16454 12980
rect 16448 12940 16896 12968
rect 16448 12928 16454 12940
rect 14277 12903 14335 12909
rect 14277 12900 14289 12903
rect 13688 12872 14289 12900
rect 13688 12860 13694 12872
rect 14277 12869 14289 12872
rect 14323 12869 14335 12903
rect 14277 12863 14335 12869
rect 14369 12903 14427 12909
rect 14369 12869 14381 12903
rect 14415 12869 14427 12903
rect 14369 12863 14427 12869
rect 15194 12860 15200 12912
rect 15252 12900 15258 12912
rect 16761 12903 16819 12909
rect 16761 12900 16773 12903
rect 15252 12872 16773 12900
rect 15252 12860 15258 12872
rect 16761 12869 16773 12872
rect 16807 12869 16819 12903
rect 16868 12900 16896 12940
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 17092 12940 17325 12968
rect 17092 12928 17098 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 17313 12931 17371 12937
rect 17865 12903 17923 12909
rect 17865 12900 17877 12903
rect 16868 12872 17877 12900
rect 16761 12863 16819 12869
rect 17865 12869 17877 12872
rect 17911 12900 17923 12903
rect 19334 12900 19340 12912
rect 17911 12872 19340 12900
rect 17911 12869 17923 12872
rect 17865 12863 17923 12869
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 9784 12804 10088 12832
rect 10152 12804 12296 12832
rect 7524 12736 8708 12764
rect 7524 12724 7530 12736
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 9784 12764 9812 12804
rect 9548 12736 9812 12764
rect 9548 12724 9554 12736
rect 9858 12724 9864 12776
rect 9916 12724 9922 12776
rect 10152 12764 10180 12804
rect 9968 12736 10180 12764
rect 5552 12668 6684 12696
rect 6932 12668 8248 12696
rect 6656 12640 6684 12668
rect 5718 12628 5724 12640
rect 4908 12600 5724 12628
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 6086 12588 6092 12640
rect 6144 12588 6150 12640
rect 6638 12588 6644 12640
rect 6696 12588 6702 12640
rect 7561 12631 7619 12637
rect 7561 12597 7573 12631
rect 7607 12628 7619 12631
rect 7926 12628 7932 12640
rect 7607 12600 7932 12628
rect 7607 12597 7619 12600
rect 7561 12591 7619 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 8076 12600 8125 12628
rect 8076 12588 8082 12600
rect 8113 12597 8125 12600
rect 8159 12597 8171 12631
rect 8220 12628 8248 12668
rect 8846 12656 8852 12708
rect 8904 12696 8910 12708
rect 9968 12696 9996 12736
rect 11698 12724 11704 12776
rect 11756 12764 11762 12776
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11756 12736 11805 12764
rect 11756 12724 11762 12736
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 12158 12724 12164 12776
rect 12216 12724 12222 12776
rect 12268 12764 12296 12804
rect 13998 12792 14004 12844
rect 14056 12792 14062 12844
rect 14094 12835 14152 12841
rect 14094 12801 14106 12835
rect 14140 12801 14152 12835
rect 14094 12795 14152 12801
rect 14507 12835 14565 12841
rect 14507 12801 14519 12835
rect 14553 12832 14565 12835
rect 14826 12832 14832 12844
rect 14553 12804 14832 12832
rect 14553 12801 14565 12804
rect 14507 12795 14565 12801
rect 12268 12736 12940 12764
rect 8904 12668 9996 12696
rect 8904 12656 8910 12668
rect 10042 12656 10048 12708
rect 10100 12696 10106 12708
rect 11146 12696 11152 12708
rect 10100 12668 11152 12696
rect 10100 12656 10106 12668
rect 11146 12656 11152 12668
rect 11204 12656 11210 12708
rect 12912 12696 12940 12736
rect 13906 12724 13912 12776
rect 13964 12764 13970 12776
rect 14109 12764 14137 12795
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 15160 12804 15485 12832
rect 15160 12792 15166 12804
rect 15473 12801 15485 12804
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 13964 12736 14137 12764
rect 13964 12724 13970 12736
rect 15010 12724 15016 12776
rect 15068 12764 15074 12776
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 15068 12736 15301 12764
rect 15068 12724 15074 12736
rect 15289 12733 15301 12736
rect 15335 12733 15347 12767
rect 15488 12764 15516 12795
rect 15838 12792 15844 12844
rect 15896 12832 15902 12844
rect 16022 12832 16028 12844
rect 15896 12804 16028 12832
rect 15896 12792 15902 12804
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16666 12832 16672 12844
rect 16132 12804 16672 12832
rect 16132 12764 16160 12804
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 17494 12792 17500 12844
rect 17552 12792 17558 12844
rect 15488 12736 16160 12764
rect 15289 12727 15347 12733
rect 16206 12724 16212 12776
rect 16264 12724 16270 12776
rect 16390 12724 16396 12776
rect 16448 12764 16454 12776
rect 17037 12767 17095 12773
rect 17037 12764 17049 12767
rect 16448 12736 17049 12764
rect 16448 12724 16454 12736
rect 17037 12733 17049 12736
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 15105 12699 15163 12705
rect 15105 12696 15117 12699
rect 12912 12668 15117 12696
rect 15105 12665 15117 12668
rect 15151 12665 15163 12699
rect 15105 12659 15163 12665
rect 15562 12656 15568 12708
rect 15620 12656 15626 12708
rect 9858 12628 9864 12640
rect 8220 12600 9864 12628
rect 8113 12591 8171 12597
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10413 12631 10471 12637
rect 10413 12597 10425 12631
rect 10459 12628 10471 12631
rect 13538 12628 13544 12640
rect 10459 12600 13544 12628
rect 10459 12597 10471 12600
rect 10413 12591 10471 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 14645 12631 14703 12637
rect 14645 12628 14657 12631
rect 13872 12600 14657 12628
rect 13872 12588 13878 12600
rect 14645 12597 14657 12600
rect 14691 12597 14703 12631
rect 14645 12591 14703 12597
rect 15286 12588 15292 12640
rect 15344 12628 15350 12640
rect 15746 12628 15752 12640
rect 15344 12600 15752 12628
rect 15344 12588 15350 12600
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 1104 12538 18860 12560
rect 1104 12486 3169 12538
rect 3221 12486 3233 12538
rect 3285 12486 3297 12538
rect 3349 12486 3361 12538
rect 3413 12486 3425 12538
rect 3477 12486 7608 12538
rect 7660 12486 7672 12538
rect 7724 12486 7736 12538
rect 7788 12486 7800 12538
rect 7852 12486 7864 12538
rect 7916 12486 12047 12538
rect 12099 12486 12111 12538
rect 12163 12486 12175 12538
rect 12227 12486 12239 12538
rect 12291 12486 12303 12538
rect 12355 12486 16486 12538
rect 16538 12486 16550 12538
rect 16602 12486 16614 12538
rect 16666 12486 16678 12538
rect 16730 12486 16742 12538
rect 16794 12486 18860 12538
rect 1104 12464 18860 12486
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 4154 12424 4160 12436
rect 3660 12396 4160 12424
rect 3660 12384 3666 12396
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 5350 12384 5356 12436
rect 5408 12384 5414 12436
rect 7742 12424 7748 12436
rect 5460 12396 7748 12424
rect 1854 12316 1860 12368
rect 1912 12356 1918 12368
rect 5460 12356 5488 12396
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 9398 12424 9404 12436
rect 8352 12396 9404 12424
rect 8352 12384 8358 12396
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 11238 12424 11244 12436
rect 9916 12396 11244 12424
rect 9916 12384 9922 12396
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 13449 12427 13507 12433
rect 13449 12424 13461 12427
rect 11848 12396 13461 12424
rect 11848 12384 11854 12396
rect 13449 12393 13461 12396
rect 13495 12424 13507 12427
rect 13906 12424 13912 12436
rect 13495 12396 13912 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 14458 12384 14464 12436
rect 14516 12424 14522 12436
rect 15654 12424 15660 12436
rect 14516 12396 15660 12424
rect 14516 12384 14522 12396
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 17405 12427 17463 12433
rect 17405 12424 17417 12427
rect 15764 12396 17417 12424
rect 1912 12328 5488 12356
rect 1912 12316 1918 12328
rect 6638 12316 6644 12368
rect 6696 12356 6702 12368
rect 7282 12356 7288 12368
rect 6696 12328 7288 12356
rect 6696 12316 6702 12328
rect 7282 12316 7288 12328
rect 7340 12316 7346 12368
rect 8312 12356 8340 12384
rect 14090 12356 14096 12368
rect 7392 12328 8340 12356
rect 10704 12328 14096 12356
rect 842 12248 848 12300
rect 900 12288 906 12300
rect 1210 12288 1216 12300
rect 900 12260 1216 12288
rect 900 12248 906 12260
rect 1210 12248 1216 12260
rect 1268 12248 1274 12300
rect 2590 12288 2596 12300
rect 2148 12260 2596 12288
rect 1118 12180 1124 12232
rect 1176 12220 1182 12232
rect 1857 12223 1915 12229
rect 1176 12192 1808 12220
rect 1176 12180 1182 12192
rect 1578 12112 1584 12164
rect 1636 12112 1642 12164
rect 1780 12152 1808 12192
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 2038 12220 2044 12232
rect 1903 12192 2044 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2148 12229 2176 12260
rect 2590 12248 2596 12260
rect 2648 12288 2654 12300
rect 3605 12291 3663 12297
rect 3605 12288 3617 12291
rect 2648 12260 3617 12288
rect 2648 12248 2654 12260
rect 3605 12257 3617 12260
rect 3651 12288 3663 12291
rect 4341 12291 4399 12297
rect 3651 12260 4292 12288
rect 3651 12257 3663 12260
rect 3605 12251 3663 12257
rect 4264 12232 4292 12260
rect 4341 12257 4353 12291
rect 4387 12288 4399 12291
rect 5077 12291 5135 12297
rect 4387 12260 4844 12288
rect 4387 12257 4399 12260
rect 4341 12251 4399 12257
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 2363 12192 2397 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2332 12152 2360 12183
rect 4246 12180 4252 12232
rect 4304 12180 4310 12232
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 2593 12155 2651 12161
rect 2593 12152 2605 12155
rect 1780 12124 2605 12152
rect 2593 12121 2605 12124
rect 2639 12121 2651 12155
rect 2593 12115 2651 12121
rect 3142 12112 3148 12164
rect 3200 12152 3206 12164
rect 4632 12152 4660 12183
rect 3200 12124 4660 12152
rect 4816 12152 4844 12260
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 5534 12288 5540 12300
rect 5123 12260 5540 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 7392 12288 7420 12328
rect 6052 12260 7420 12288
rect 6052 12248 6058 12260
rect 7742 12248 7748 12300
rect 7800 12288 7806 12300
rect 8389 12291 8447 12297
rect 7800 12260 8064 12288
rect 7800 12248 7806 12260
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5350 12220 5356 12232
rect 4939 12192 5356 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 8036 12229 8064 12260
rect 8389 12257 8401 12291
rect 8435 12288 8447 12291
rect 10704 12288 10732 12328
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 8435 12260 10732 12288
rect 10781 12291 10839 12297
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 11698 12288 11704 12300
rect 10827 12260 11704 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11698 12248 11704 12260
rect 11756 12288 11762 12300
rect 12618 12288 12624 12300
rect 11756 12260 12624 12288
rect 11756 12248 11762 12260
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 15764 12288 15792 12396
rect 17405 12393 17417 12396
rect 17451 12393 17463 12427
rect 17405 12387 17463 12393
rect 13964 12260 15792 12288
rect 13964 12248 13970 12260
rect 15930 12248 15936 12300
rect 15988 12248 15994 12300
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7064 12192 7849 12220
rect 7064 12180 7070 12192
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9227 12220 9352 12222
rect 9490 12220 9496 12232
rect 9180 12194 9496 12220
rect 9180 12192 9255 12194
rect 9324 12192 9496 12194
rect 9180 12180 9186 12192
rect 9490 12180 9496 12192
rect 9548 12180 9554 12232
rect 11054 12180 11060 12232
rect 11112 12180 11118 12232
rect 11790 12180 11796 12232
rect 11848 12180 11854 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 14826 12220 14832 12232
rect 14415 12192 14832 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15654 12180 15660 12232
rect 15712 12180 15718 12232
rect 5810 12152 5816 12164
rect 4816 12124 5816 12152
rect 3200 12112 3206 12124
rect 5810 12112 5816 12124
rect 5868 12112 5874 12164
rect 7190 12112 7196 12164
rect 7248 12152 7254 12164
rect 7466 12152 7472 12164
rect 7248 12124 7472 12152
rect 7248 12112 7254 12124
rect 7466 12112 7472 12124
rect 7524 12112 7530 12164
rect 7742 12112 7748 12164
rect 7800 12112 7806 12164
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 8478 12152 8484 12164
rect 8168 12124 8484 12152
rect 8168 12112 8174 12124
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 10505 12155 10563 12161
rect 10505 12121 10517 12155
rect 10551 12152 10563 12155
rect 13262 12152 13268 12164
rect 10551 12124 13268 12152
rect 10551 12121 10563 12124
rect 10505 12115 10563 12121
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 15470 12152 15476 12164
rect 13740 12124 15476 12152
rect 1670 12044 1676 12096
rect 1728 12084 1734 12096
rect 1949 12087 2007 12093
rect 1949 12084 1961 12087
rect 1728 12056 1961 12084
rect 1728 12044 1734 12056
rect 1949 12053 1961 12056
rect 1995 12053 2007 12087
rect 1949 12047 2007 12053
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 3053 12087 3111 12093
rect 3053 12084 3065 12087
rect 2924 12056 3065 12084
rect 2924 12044 2930 12056
rect 3053 12053 3065 12056
rect 3099 12084 3111 12087
rect 4338 12084 4344 12096
rect 3099 12056 4344 12084
rect 3099 12053 3111 12056
rect 3053 12047 3111 12053
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 5077 12087 5135 12093
rect 5077 12053 5089 12087
rect 5123 12084 5135 12087
rect 5166 12084 5172 12096
rect 5123 12056 5172 12084
rect 5123 12053 5135 12056
rect 5077 12047 5135 12053
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 5721 12087 5779 12093
rect 5721 12053 5733 12087
rect 5767 12084 5779 12087
rect 6270 12084 6276 12096
rect 5767 12056 6276 12084
rect 5767 12053 5779 12056
rect 5721 12047 5779 12053
rect 6270 12044 6276 12056
rect 6328 12084 6334 12096
rect 6457 12087 6515 12093
rect 6457 12084 6469 12087
rect 6328 12056 6469 12084
rect 6328 12044 6334 12056
rect 6457 12053 6469 12056
rect 6503 12084 6515 12087
rect 6546 12084 6552 12096
rect 6503 12056 6552 12084
rect 6503 12053 6515 12056
rect 6457 12047 6515 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 8297 12087 8355 12093
rect 8297 12053 8309 12087
rect 8343 12084 8355 12087
rect 8754 12084 8760 12096
rect 8343 12056 8760 12084
rect 8343 12053 8355 12056
rect 8297 12047 8355 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 9033 12087 9091 12093
rect 9033 12053 9045 12087
rect 9079 12084 9091 12087
rect 9582 12084 9588 12096
rect 9079 12056 9588 12084
rect 9079 12053 9091 12056
rect 9033 12047 9091 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 10965 12087 11023 12093
rect 10965 12084 10977 12087
rect 10468 12056 10977 12084
rect 10468 12044 10474 12056
rect 10965 12053 10977 12056
rect 11011 12053 11023 12087
rect 10965 12047 11023 12053
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11698 12084 11704 12096
rect 11112 12056 11704 12084
rect 11112 12044 11118 12056
rect 11698 12044 11704 12056
rect 11756 12084 11762 12096
rect 13740 12084 13768 12124
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 16040 12124 16422 12152
rect 11756 12056 13768 12084
rect 13909 12087 13967 12093
rect 11756 12044 11762 12056
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14182 12084 14188 12096
rect 13955 12056 14188 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14516 12056 14657 12084
rect 14516 12044 14522 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15381 12087 15439 12093
rect 15381 12084 15393 12087
rect 15344 12056 15393 12084
rect 15344 12044 15350 12056
rect 15381 12053 15393 12056
rect 15427 12084 15439 12087
rect 16040 12084 16068 12124
rect 15427 12056 16068 12084
rect 15427 12053 15439 12056
rect 15381 12047 15439 12053
rect 1104 11994 18860 12016
rect 1104 11942 3829 11994
rect 3881 11942 3893 11994
rect 3945 11942 3957 11994
rect 4009 11942 4021 11994
rect 4073 11942 4085 11994
rect 4137 11942 8268 11994
rect 8320 11942 8332 11994
rect 8384 11942 8396 11994
rect 8448 11942 8460 11994
rect 8512 11942 8524 11994
rect 8576 11942 12707 11994
rect 12759 11942 12771 11994
rect 12823 11942 12835 11994
rect 12887 11942 12899 11994
rect 12951 11942 12963 11994
rect 13015 11942 17146 11994
rect 17198 11942 17210 11994
rect 17262 11942 17274 11994
rect 17326 11942 17338 11994
rect 17390 11942 17402 11994
rect 17454 11942 18860 11994
rect 1104 11920 18860 11942
rect 566 11840 572 11892
rect 624 11880 630 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 624 11852 6469 11880
rect 624 11840 630 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 7098 11880 7104 11892
rect 6457 11843 6515 11849
rect 6564 11852 7104 11880
rect 2593 11815 2651 11821
rect 2593 11781 2605 11815
rect 2639 11812 2651 11815
rect 2866 11812 2872 11824
rect 2639 11784 2872 11812
rect 2639 11781 2651 11784
rect 2593 11775 2651 11781
rect 2866 11772 2872 11784
rect 2924 11772 2930 11824
rect 3329 11815 3387 11821
rect 3329 11781 3341 11815
rect 3375 11812 3387 11815
rect 3694 11812 3700 11824
rect 3375 11784 3700 11812
rect 3375 11781 3387 11784
rect 3329 11775 3387 11781
rect 1670 11704 1676 11756
rect 1728 11704 1734 11756
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11744 1823 11747
rect 2130 11744 2136 11756
rect 1811 11716 2136 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 2406 11753 2412 11756
rect 2404 11744 2412 11753
rect 2367 11716 2412 11744
rect 2404 11707 2412 11716
rect 2406 11704 2412 11707
rect 2464 11704 2470 11756
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 2041 11679 2099 11685
rect 2041 11676 2053 11679
rect 2004 11648 2053 11676
rect 2004 11636 2010 11648
rect 2041 11645 2053 11648
rect 2087 11645 2099 11679
rect 2516 11676 2544 11707
rect 2774 11704 2780 11756
rect 2832 11704 2838 11756
rect 3344 11676 3372 11775
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 4062 11772 4068 11824
rect 4120 11772 4126 11824
rect 3970 11704 3976 11756
rect 4028 11704 4034 11756
rect 4080 11744 4108 11772
rect 4080 11716 4200 11744
rect 4172 11685 4200 11716
rect 4614 11704 4620 11756
rect 4672 11744 4678 11756
rect 5350 11744 5356 11756
rect 4672 11716 5356 11744
rect 4672 11704 4678 11716
rect 5350 11704 5356 11716
rect 5408 11744 5414 11756
rect 6564 11753 6592 11852
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7926 11840 7932 11892
rect 7984 11840 7990 11892
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 9214 11880 9220 11892
rect 8076 11852 9220 11880
rect 8076 11840 8082 11852
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9398 11840 9404 11892
rect 9456 11880 9462 11892
rect 13906 11880 13912 11892
rect 9456 11852 13912 11880
rect 9456 11840 9462 11852
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 16390 11880 16396 11892
rect 15528 11852 16396 11880
rect 15528 11840 15534 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 16761 11883 16819 11889
rect 16761 11849 16773 11883
rect 16807 11880 16819 11883
rect 16850 11880 16856 11892
rect 16807 11852 16856 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 8846 11812 8852 11824
rect 6656 11784 6961 11812
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 5408 11716 6561 11744
rect 5408 11704 5414 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 2516 11648 3372 11676
rect 4065 11679 4123 11685
rect 2041 11639 2099 11645
rect 4065 11645 4077 11679
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 5534 11676 5540 11688
rect 5491 11648 5540 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 1489 11611 1547 11617
rect 1489 11577 1501 11611
rect 1535 11608 1547 11611
rect 2498 11608 2504 11620
rect 1535 11580 2504 11608
rect 1535 11577 1547 11580
rect 1489 11571 1547 11577
rect 2498 11568 2504 11580
rect 2556 11568 2562 11620
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 3605 11611 3663 11617
rect 3605 11608 3617 11611
rect 2832 11580 3617 11608
rect 2832 11568 2838 11580
rect 3605 11577 3617 11580
rect 3651 11577 3663 11611
rect 3605 11571 3663 11577
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 1854 11540 1860 11552
rect 1636 11512 1860 11540
rect 1636 11500 1642 11512
rect 1854 11500 1860 11512
rect 1912 11540 1918 11552
rect 1949 11543 2007 11549
rect 1949 11540 1961 11543
rect 1912 11512 1961 11540
rect 1912 11500 1918 11512
rect 1949 11509 1961 11512
rect 1995 11509 2007 11543
rect 1949 11503 2007 11509
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 3142 11540 3148 11552
rect 2271 11512 3148 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 4080 11540 4108 11639
rect 5534 11636 5540 11648
rect 5592 11676 5598 11688
rect 6656 11676 6684 11784
rect 6822 11704 6828 11756
rect 6880 11704 6886 11756
rect 6933 11753 6961 11784
rect 7116 11784 8852 11812
rect 7116 11753 7144 11784
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 11330 11772 11336 11824
rect 11388 11812 11394 11824
rect 14093 11815 14151 11821
rect 14093 11812 14105 11815
rect 11388 11784 14105 11812
rect 11388 11772 11394 11784
rect 14093 11781 14105 11784
rect 14139 11781 14151 11815
rect 14093 11775 14151 11781
rect 16209 11815 16267 11821
rect 16209 11781 16221 11815
rect 16255 11812 16267 11815
rect 16298 11812 16304 11824
rect 16255 11784 16304 11812
rect 16255 11781 16267 11784
rect 16209 11775 16267 11781
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 16482 11772 16488 11824
rect 16540 11772 16546 11824
rect 17310 11812 17316 11824
rect 16776 11784 17316 11812
rect 6918 11747 6976 11753
rect 6918 11713 6930 11747
rect 6964 11713 6976 11747
rect 6918 11707 6976 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11744 7619 11747
rect 9214 11744 9220 11756
rect 7607 11716 9220 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 9214 11704 9220 11716
rect 9272 11744 9278 11756
rect 10962 11744 10968 11756
rect 9272 11716 10968 11744
rect 9272 11704 9278 11716
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11790 11704 11796 11756
rect 11848 11704 11854 11756
rect 13722 11744 13728 11756
rect 13280 11716 13728 11744
rect 5592 11648 6684 11676
rect 6733 11679 6791 11685
rect 5592 11636 5598 11648
rect 6733 11645 6745 11679
rect 6779 11676 6791 11679
rect 6779 11648 7031 11676
rect 6779 11645 6791 11648
rect 6733 11639 6791 11645
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 5258 11608 5264 11620
rect 4764 11580 5264 11608
rect 4764 11568 4770 11580
rect 5258 11568 5264 11580
rect 5316 11608 5322 11620
rect 7003 11608 7031 11648
rect 7282 11636 7288 11688
rect 7340 11636 7346 11688
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11676 7527 11679
rect 7650 11676 7656 11688
rect 7515 11648 7656 11676
rect 7515 11645 7527 11648
rect 7469 11639 7527 11645
rect 7650 11636 7656 11648
rect 7708 11676 7714 11688
rect 8386 11676 8392 11688
rect 7708 11648 8392 11676
rect 7708 11636 7714 11648
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8570 11636 8576 11688
rect 8628 11676 8634 11688
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 8628 11648 10701 11676
rect 8628 11636 8634 11648
rect 10689 11645 10701 11648
rect 10735 11676 10747 11679
rect 11808 11676 11836 11704
rect 10735 11648 11836 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 13078 11636 13084 11688
rect 13136 11676 13142 11688
rect 13280 11685 13308 11716
rect 13722 11704 13728 11716
rect 13780 11744 13786 11756
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13780 11716 13921 11744
rect 13780 11704 13786 11716
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 13909 11707 13967 11713
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14734 11744 14740 11756
rect 14240 11716 14740 11744
rect 14240 11704 14246 11716
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16500 11744 16528 11772
rect 16776 11753 16804 11784
rect 17310 11772 17316 11784
rect 17368 11772 17374 11824
rect 16163 11716 16528 11744
rect 16761 11747 16819 11753
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16761 11713 16773 11747
rect 16807 11713 16819 11747
rect 16761 11707 16819 11713
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 17000 11716 17693 11744
rect 17000 11704 17006 11716
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 13136 11648 13277 11676
rect 13136 11636 13142 11648
rect 13265 11645 13277 11648
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11645 13507 11679
rect 13449 11639 13507 11645
rect 11054 11608 11060 11620
rect 5316 11580 6960 11608
rect 7003 11580 11060 11608
rect 5316 11568 5322 11580
rect 4890 11540 4896 11552
rect 4080 11512 4896 11540
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5350 11500 5356 11552
rect 5408 11540 5414 11552
rect 5721 11543 5779 11549
rect 5721 11540 5733 11543
rect 5408 11512 5733 11540
rect 5408 11500 5414 11512
rect 5721 11509 5733 11512
rect 5767 11509 5779 11543
rect 5721 11503 5779 11509
rect 6086 11500 6092 11552
rect 6144 11540 6150 11552
rect 6181 11543 6239 11549
rect 6181 11540 6193 11543
rect 6144 11512 6193 11540
rect 6144 11500 6150 11512
rect 6181 11509 6193 11512
rect 6227 11540 6239 11543
rect 6822 11540 6828 11552
rect 6227 11512 6828 11540
rect 6227 11509 6239 11512
rect 6181 11503 6239 11509
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 6932 11540 6960 11580
rect 11054 11568 11060 11580
rect 11112 11568 11118 11620
rect 12894 11608 12900 11620
rect 11256 11580 12900 11608
rect 8570 11540 8576 11552
rect 6932 11512 8576 11540
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 8849 11543 8907 11549
rect 8849 11509 8861 11543
rect 8895 11540 8907 11543
rect 9214 11540 9220 11552
rect 8895 11512 9220 11540
rect 8895 11509 8907 11512
rect 8849 11503 8907 11509
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 11256 11540 11284 11580
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 13464 11608 13492 11639
rect 14458 11636 14464 11688
rect 14516 11676 14522 11688
rect 15841 11679 15899 11685
rect 15841 11676 15853 11679
rect 14516 11648 15853 11676
rect 14516 11636 14522 11648
rect 15841 11645 15853 11648
rect 15887 11645 15899 11679
rect 15841 11639 15899 11645
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 16485 11679 16543 11685
rect 16485 11645 16497 11679
rect 16531 11676 16543 11679
rect 18138 11676 18144 11688
rect 16531 11648 18144 11676
rect 16531 11645 16543 11648
rect 16485 11639 16543 11645
rect 13004 11580 14872 11608
rect 9364 11512 11284 11540
rect 9364 11500 9370 11512
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 13004 11549 13032 11580
rect 12989 11543 13047 11549
rect 12989 11540 13001 11543
rect 11388 11512 13001 11540
rect 11388 11500 11394 11512
rect 12989 11509 13001 11512
rect 13035 11509 13047 11543
rect 12989 11503 13047 11509
rect 13630 11500 13636 11552
rect 13688 11500 13694 11552
rect 14844 11540 14872 11580
rect 16022 11540 16028 11552
rect 14844 11512 16028 11540
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 16224 11540 16252 11639
rect 16408 11608 16436 11639
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 17494 11608 17500 11620
rect 16408 11580 17500 11608
rect 17494 11568 17500 11580
rect 17552 11568 17558 11620
rect 17313 11543 17371 11549
rect 17313 11540 17325 11543
rect 16224 11512 17325 11540
rect 17313 11509 17325 11512
rect 17359 11540 17371 11543
rect 18414 11540 18420 11552
rect 17359 11512 18420 11540
rect 17359 11509 17371 11512
rect 17313 11503 17371 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 1104 11450 18860 11472
rect 1104 11398 3169 11450
rect 3221 11398 3233 11450
rect 3285 11398 3297 11450
rect 3349 11398 3361 11450
rect 3413 11398 3425 11450
rect 3477 11398 7608 11450
rect 7660 11398 7672 11450
rect 7724 11398 7736 11450
rect 7788 11398 7800 11450
rect 7852 11398 7864 11450
rect 7916 11398 12047 11450
rect 12099 11398 12111 11450
rect 12163 11398 12175 11450
rect 12227 11398 12239 11450
rect 12291 11398 12303 11450
rect 12355 11398 16486 11450
rect 16538 11398 16550 11450
rect 16602 11398 16614 11450
rect 16666 11398 16678 11450
rect 16730 11398 16742 11450
rect 16794 11398 18860 11450
rect 1104 11376 18860 11398
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11336 4399 11339
rect 4614 11336 4620 11348
rect 4387 11308 4620 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6822 11336 6828 11348
rect 5868 11308 6828 11336
rect 5868 11296 5874 11308
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 7558 11336 7564 11348
rect 7340 11308 7564 11336
rect 7340 11296 7346 11308
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 8404 11308 9137 11336
rect 1302 11228 1308 11280
rect 1360 11268 1366 11280
rect 1581 11271 1639 11277
rect 1581 11268 1593 11271
rect 1360 11240 1593 11268
rect 1360 11228 1366 11240
rect 1581 11237 1593 11240
rect 1627 11237 1639 11271
rect 1581 11231 1639 11237
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4709 11271 4767 11277
rect 4709 11268 4721 11271
rect 4028 11240 4721 11268
rect 4028 11228 4034 11240
rect 4709 11237 4721 11240
rect 4755 11268 4767 11271
rect 5994 11268 6000 11280
rect 4755 11240 6000 11268
rect 4755 11237 4767 11240
rect 4709 11231 4767 11237
rect 5994 11228 6000 11240
rect 6052 11268 6058 11280
rect 6270 11268 6276 11280
rect 6052 11240 6276 11268
rect 6052 11228 6058 11240
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 8404 11268 8432 11308
rect 9125 11305 9137 11308
rect 9171 11336 9183 11339
rect 11330 11336 11336 11348
rect 9171 11308 11336 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11425 11339 11483 11345
rect 11425 11305 11437 11339
rect 11471 11336 11483 11339
rect 11514 11336 11520 11348
rect 11471 11308 11520 11336
rect 11471 11305 11483 11308
rect 11425 11299 11483 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 15010 11296 15016 11348
rect 15068 11336 15074 11348
rect 15197 11339 15255 11345
rect 15197 11336 15209 11339
rect 15068 11308 15209 11336
rect 15068 11296 15074 11308
rect 15197 11305 15209 11308
rect 15243 11336 15255 11339
rect 15286 11336 15292 11348
rect 15243 11308 15292 11336
rect 15243 11305 15255 11308
rect 15197 11299 15255 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15930 11296 15936 11348
rect 15988 11296 15994 11348
rect 8128 11240 8432 11268
rect 2590 11160 2596 11212
rect 2648 11200 2654 11212
rect 3329 11203 3387 11209
rect 3329 11200 3341 11203
rect 2648 11172 3341 11200
rect 2648 11160 2654 11172
rect 3329 11169 3341 11172
rect 3375 11169 3387 11203
rect 3329 11163 3387 11169
rect 3605 11203 3663 11209
rect 3605 11169 3617 11203
rect 3651 11200 3663 11203
rect 4154 11200 4160 11212
rect 3651 11172 4160 11200
rect 3651 11169 3663 11172
rect 3605 11163 3663 11169
rect 4154 11160 4160 11172
rect 4212 11200 4218 11212
rect 6546 11200 6552 11212
rect 4212 11172 6552 11200
rect 4212 11160 4218 11172
rect 6546 11160 6552 11172
rect 6604 11200 6610 11212
rect 7554 11203 7612 11209
rect 7554 11200 7566 11203
rect 6604 11172 7566 11200
rect 6604 11160 6610 11172
rect 7554 11169 7566 11172
rect 7600 11169 7612 11203
rect 8128 11200 8156 11240
rect 9030 11228 9036 11280
rect 9088 11228 9094 11280
rect 9398 11228 9404 11280
rect 9456 11268 9462 11280
rect 9456 11240 14320 11268
rect 9456 11228 9462 11240
rect 9048 11200 9076 11228
rect 7554 11163 7612 11169
rect 7668 11172 8156 11200
rect 8496 11172 9076 11200
rect 7668 11144 7696 11172
rect 1394 11092 1400 11144
rect 1452 11132 1458 11144
rect 2038 11132 2044 11144
rect 1452 11104 2044 11132
rect 1452 11092 1458 11104
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 5994 11132 6000 11144
rect 4580 11104 6000 11132
rect 4580 11092 4586 11104
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 7650 11092 7656 11144
rect 7708 11092 7714 11144
rect 7834 11092 7840 11144
rect 7892 11092 7898 11144
rect 8110 11092 8116 11144
rect 8168 11092 8174 11144
rect 8309 11135 8367 11141
rect 8309 11101 8321 11135
rect 8355 11132 8367 11135
rect 8496 11132 8524 11172
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 13722 11200 13728 11212
rect 9548 11172 13728 11200
rect 9548 11160 9554 11172
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 8355 11104 8524 11132
rect 8665 11135 8723 11141
rect 8355 11101 8367 11104
rect 8309 11095 8367 11101
rect 8665 11101 8677 11135
rect 8711 11132 8723 11135
rect 9306 11132 9312 11144
rect 8711 11104 9312 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 1670 11024 1676 11076
rect 1728 11064 1734 11076
rect 1946 11064 1952 11076
rect 1728 11036 1952 11064
rect 1728 11024 1734 11036
rect 1946 11024 1952 11036
rect 2004 11024 2010 11076
rect 2682 11024 2688 11076
rect 2740 11024 2746 11076
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 5353 11067 5411 11073
rect 5353 11064 5365 11067
rect 5316 11036 5365 11064
rect 5316 11024 5322 11036
rect 5353 11033 5365 11036
rect 5399 11033 5411 11067
rect 5353 11027 5411 11033
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 5776 11036 6118 11064
rect 5776 11024 5782 11036
rect 7282 11024 7288 11076
rect 7340 11024 7346 11076
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 8680 11064 8708 11095
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 12158 11132 12164 11144
rect 9824 11104 12164 11132
rect 9824 11092 9830 11104
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 12897 11135 12955 11141
rect 12897 11132 12909 11135
rect 12676 11104 12909 11132
rect 12676 11092 12682 11104
rect 12897 11101 12909 11104
rect 12943 11101 12955 11135
rect 12897 11095 12955 11101
rect 13630 11092 13636 11144
rect 13688 11132 13694 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13688 11104 14197 11132
rect 13688 11092 13694 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14292 11132 14320 11240
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 15028 11200 15056 11296
rect 16022 11228 16028 11280
rect 16080 11268 16086 11280
rect 16666 11268 16672 11280
rect 16080 11240 16672 11268
rect 16080 11228 16086 11240
rect 16666 11228 16672 11240
rect 16724 11228 16730 11280
rect 16945 11271 17003 11277
rect 16945 11237 16957 11271
rect 16991 11268 17003 11271
rect 17862 11268 17868 11280
rect 16991 11240 17868 11268
rect 16991 11237 17003 11240
rect 16945 11231 17003 11237
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 14507 11172 15056 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 14350 11135 14408 11141
rect 14350 11132 14362 11135
rect 14292 11104 14362 11132
rect 14185 11095 14243 11101
rect 14350 11101 14362 11104
rect 14396 11132 14408 11135
rect 14396 11104 14504 11132
rect 14396 11101 14408 11104
rect 14350 11095 14408 11101
rect 7616 11036 8708 11064
rect 7616 11024 7622 11036
rect 9582 11024 9588 11076
rect 9640 11064 9646 11076
rect 13446 11064 13452 11076
rect 9640 11036 13452 11064
rect 9640 11024 9646 11036
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 13541 11067 13599 11073
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 13587 11036 13676 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 1854 10956 1860 11008
rect 1912 10956 1918 11008
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 4062 10996 4068 11008
rect 3476 10968 4068 10996
rect 3476 10956 3482 10968
rect 4062 10956 4068 10968
rect 4120 10996 4126 11008
rect 5077 10999 5135 11005
rect 5077 10996 5089 10999
rect 4120 10968 5089 10996
rect 4120 10956 4126 10968
rect 5077 10965 5089 10968
rect 5123 10996 5135 10999
rect 6546 10996 6552 11008
rect 5123 10968 6552 10996
rect 5123 10965 5135 10968
rect 5077 10959 5135 10965
rect 6546 10956 6552 10968
rect 6604 10996 6610 11008
rect 7576 10996 7604 11024
rect 6604 10968 7604 10996
rect 6604 10956 6610 10968
rect 7926 10956 7932 11008
rect 7984 10996 7990 11008
rect 8021 10999 8079 11005
rect 8021 10996 8033 10999
rect 7984 10968 8033 10996
rect 7984 10956 7990 10968
rect 8021 10965 8033 10968
rect 8067 10965 8079 10999
rect 8021 10959 8079 10965
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 11054 10996 11060 11008
rect 8168 10968 11060 10996
rect 8168 10956 8174 10968
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 13648 10996 13676 11036
rect 13722 11024 13728 11076
rect 13780 11024 13786 11076
rect 14476 11064 14504 11104
rect 14550 11092 14556 11144
rect 14608 11092 14614 11144
rect 14642 11092 14648 11144
rect 14700 11132 14706 11144
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 14700 11104 14749 11132
rect 14700 11092 14706 11104
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 14918 11092 14924 11144
rect 14976 11092 14982 11144
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 16390 11132 16396 11144
rect 16347 11104 16396 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11101 16543 11135
rect 16485 11095 16543 11101
rect 15565 11067 15623 11073
rect 15565 11064 15577 11067
rect 14476 11036 15577 11064
rect 15565 11033 15577 11036
rect 15611 11064 15623 11067
rect 15746 11064 15752 11076
rect 15611 11036 15752 11064
rect 15611 11033 15623 11036
rect 15565 11027 15623 11033
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 16500 11064 16528 11095
rect 16574 11092 16580 11144
rect 16632 11092 16638 11144
rect 16703 11135 16761 11141
rect 16703 11101 16715 11135
rect 16749 11132 16761 11135
rect 16942 11132 16948 11144
rect 16749 11104 16948 11132
rect 16749 11101 16761 11104
rect 16703 11095 16761 11101
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17681 11135 17739 11141
rect 17681 11101 17693 11135
rect 17727 11132 17739 11135
rect 18414 11132 18420 11144
rect 17727 11104 18420 11132
rect 17727 11101 17739 11104
rect 17681 11095 17739 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 16132 11036 16528 11064
rect 16132 11008 16160 11036
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17862 11064 17868 11076
rect 17368 11036 17868 11064
rect 17368 11024 17374 11036
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 13906 10996 13912 11008
rect 13648 10968 13912 10996
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 15194 10996 15200 11008
rect 14884 10968 15200 10996
rect 14884 10956 14890 10968
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 16114 10956 16120 11008
rect 16172 10956 16178 11008
rect 1104 10906 18860 10928
rect 1104 10854 3829 10906
rect 3881 10854 3893 10906
rect 3945 10854 3957 10906
rect 4009 10854 4021 10906
rect 4073 10854 4085 10906
rect 4137 10854 8268 10906
rect 8320 10854 8332 10906
rect 8384 10854 8396 10906
rect 8448 10854 8460 10906
rect 8512 10854 8524 10906
rect 8576 10854 12707 10906
rect 12759 10854 12771 10906
rect 12823 10854 12835 10906
rect 12887 10854 12899 10906
rect 12951 10854 12963 10906
rect 13015 10854 17146 10906
rect 17198 10854 17210 10906
rect 17262 10854 17274 10906
rect 17326 10854 17338 10906
rect 17390 10854 17402 10906
rect 17454 10854 18860 10906
rect 1104 10832 18860 10854
rect 1857 10795 1915 10801
rect 1857 10761 1869 10795
rect 1903 10792 1915 10795
rect 2222 10792 2228 10804
rect 1903 10764 2228 10792
rect 1903 10761 1915 10764
rect 1857 10755 1915 10761
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2869 10795 2927 10801
rect 2869 10792 2881 10795
rect 2464 10764 2881 10792
rect 2464 10752 2470 10764
rect 2869 10761 2881 10764
rect 2915 10792 2927 10795
rect 3326 10792 3332 10804
rect 2915 10764 3332 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 3697 10795 3755 10801
rect 3697 10761 3709 10795
rect 3743 10792 3755 10795
rect 4614 10792 4620 10804
rect 3743 10764 4620 10792
rect 3743 10761 3755 10764
rect 3697 10755 3755 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 5258 10792 5264 10804
rect 4856 10764 5264 10792
rect 4856 10752 4862 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 6454 10792 6460 10804
rect 5500 10764 6460 10792
rect 5500 10752 5506 10764
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 6696 10764 7297 10792
rect 6696 10752 6702 10764
rect 7285 10761 7297 10764
rect 7331 10792 7343 10795
rect 7466 10792 7472 10804
rect 7331 10764 7472 10792
rect 7331 10761 7343 10764
rect 7285 10755 7343 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 9398 10792 9404 10804
rect 7800 10764 9404 10792
rect 7800 10752 7806 10764
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 9582 10792 9588 10804
rect 9508 10764 9588 10792
rect 1578 10684 1584 10736
rect 1636 10724 1642 10736
rect 1946 10724 1952 10736
rect 1636 10696 1952 10724
rect 1636 10684 1642 10696
rect 1946 10684 1952 10696
rect 2004 10724 2010 10736
rect 2501 10727 2559 10733
rect 2501 10724 2513 10727
rect 2004 10696 2513 10724
rect 2004 10684 2010 10696
rect 2501 10693 2513 10696
rect 2547 10693 2559 10727
rect 2501 10687 2559 10693
rect 3605 10727 3663 10733
rect 3605 10693 3617 10727
rect 3651 10724 3663 10727
rect 4816 10724 4844 10752
rect 5718 10724 5724 10736
rect 3651 10696 4844 10724
rect 5658 10696 5724 10724
rect 3651 10693 3663 10696
rect 3605 10687 3663 10693
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 6362 10684 6368 10736
rect 6420 10724 6426 10736
rect 7098 10724 7104 10736
rect 6420 10696 7104 10724
rect 6420 10684 6426 10696
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 7650 10724 7656 10736
rect 7432 10696 7656 10724
rect 7432 10684 7438 10696
rect 7650 10684 7656 10696
rect 7708 10684 7714 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 8202 10724 8208 10736
rect 7892 10696 8208 10724
rect 7892 10684 7898 10696
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 9508 10724 9536 10764
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 10597 10795 10655 10801
rect 10597 10761 10609 10795
rect 10643 10792 10655 10795
rect 10778 10792 10784 10804
rect 10643 10764 10784 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 10612 10724 10640 10755
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11977 10795 12035 10801
rect 11977 10792 11989 10795
rect 11296 10764 11989 10792
rect 11296 10752 11302 10764
rect 11977 10761 11989 10764
rect 12023 10761 12035 10795
rect 11977 10755 12035 10761
rect 12618 10752 12624 10804
rect 12676 10792 12682 10804
rect 13538 10792 13544 10804
rect 12676 10764 13544 10792
rect 12676 10752 12682 10764
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 16816 10764 18061 10792
rect 16816 10752 16822 10764
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 8307 10696 8703 10724
rect 1394 10616 1400 10668
rect 1452 10616 1458 10668
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2866 10656 2872 10668
rect 2271 10628 2872 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 6181 10659 6239 10665
rect 6181 10625 6193 10659
rect 6227 10656 6239 10659
rect 6730 10656 6736 10668
rect 6227 10628 6736 10656
rect 6227 10625 6239 10628
rect 6181 10619 6239 10625
rect 6730 10616 6736 10628
rect 6788 10656 6794 10668
rect 8307 10656 8335 10696
rect 6788 10628 8335 10656
rect 6788 10616 6794 10628
rect 8570 10616 8576 10668
rect 8628 10616 8634 10668
rect 2130 10548 2136 10600
rect 2188 10548 2194 10600
rect 3418 10548 3424 10600
rect 3476 10588 3482 10600
rect 3970 10588 3976 10600
rect 3476 10560 3976 10588
rect 3476 10548 3482 10560
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10588 4491 10591
rect 5166 10588 5172 10600
rect 4479 10560 5172 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 8675 10588 8703 10696
rect 9140 10696 9536 10724
rect 9600 10696 10640 10724
rect 9140 10665 9168 10696
rect 9600 10668 9628 10696
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 11882 10724 11888 10736
rect 11388 10696 11888 10724
rect 11388 10684 11394 10696
rect 11882 10684 11888 10696
rect 11940 10684 11946 10736
rect 14550 10724 14556 10736
rect 11992 10696 14556 10724
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 9582 10656 9588 10668
rect 9447 10628 9588 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 9674 10616 9680 10668
rect 9732 10616 9738 10668
rect 11992 10656 12020 10696
rect 14550 10684 14556 10696
rect 14608 10684 14614 10736
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 14921 10727 14979 10733
rect 14921 10724 14933 10727
rect 14700 10696 14933 10724
rect 14700 10684 14706 10696
rect 14921 10693 14933 10696
rect 14967 10724 14979 10727
rect 17586 10724 17592 10736
rect 14967 10696 17592 10724
rect 14967 10693 14979 10696
rect 14921 10687 14979 10693
rect 17586 10684 17592 10696
rect 17644 10724 17650 10736
rect 18874 10724 18880 10736
rect 17644 10696 18880 10724
rect 17644 10684 17650 10696
rect 18874 10684 18880 10696
rect 18932 10684 18938 10736
rect 10152 10628 12020 10656
rect 10152 10588 10180 10628
rect 12802 10616 12808 10668
rect 12860 10616 12866 10668
rect 13538 10616 13544 10668
rect 13596 10656 13602 10668
rect 14461 10659 14519 10665
rect 14461 10656 14473 10659
rect 13596 10628 14473 10656
rect 13596 10616 13602 10628
rect 14461 10625 14473 10628
rect 14507 10656 14519 10659
rect 16482 10656 16488 10668
rect 14507 10628 16488 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16666 10616 16672 10668
rect 16724 10656 16730 10668
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16724 10628 16865 10656
rect 16724 10616 16730 10628
rect 16853 10625 16865 10628
rect 16899 10656 16911 10659
rect 17402 10656 17408 10668
rect 16899 10628 17408 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 17954 10616 17960 10668
rect 18012 10616 18018 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 18414 10656 18420 10668
rect 18371 10628 18420 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 7156 10560 8616 10588
rect 8675 10560 10180 10588
rect 7156 10548 7162 10560
rect 1578 10480 1584 10532
rect 1636 10480 1642 10532
rect 4062 10480 4068 10532
rect 4120 10480 4126 10532
rect 7469 10523 7527 10529
rect 5828 10492 7420 10520
rect 2225 10455 2283 10461
rect 2225 10421 2237 10455
rect 2271 10452 2283 10455
rect 2314 10452 2320 10464
rect 2271 10424 2320 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 5828 10452 5856 10492
rect 2924 10424 5856 10452
rect 2924 10412 2930 10424
rect 5902 10412 5908 10464
rect 5960 10452 5966 10464
rect 7098 10452 7104 10464
rect 5960 10424 7104 10452
rect 5960 10412 5966 10424
rect 7098 10412 7104 10424
rect 7156 10452 7162 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 7156 10424 7297 10452
rect 7156 10412 7162 10424
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 7392 10452 7420 10492
rect 7469 10489 7481 10523
rect 7515 10520 7527 10523
rect 7515 10492 8432 10520
rect 7515 10489 7527 10492
rect 7469 10483 7527 10489
rect 7650 10452 7656 10464
rect 7392 10424 7656 10452
rect 7285 10415 7343 10421
rect 7650 10412 7656 10424
rect 7708 10452 7714 10464
rect 8110 10452 8116 10464
rect 7708 10424 8116 10452
rect 7708 10412 7714 10424
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8202 10412 8208 10464
rect 8260 10412 8266 10464
rect 8404 10452 8432 10492
rect 8478 10480 8484 10532
rect 8536 10480 8542 10532
rect 8588 10520 8616 10560
rect 10226 10548 10232 10600
rect 10284 10548 10290 10600
rect 11514 10548 11520 10600
rect 11572 10588 11578 10600
rect 11974 10588 11980 10600
rect 11572 10560 11980 10588
rect 11572 10548 11578 10560
rect 11974 10548 11980 10560
rect 12032 10588 12038 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 12032 10560 12081 10588
rect 12032 10548 12038 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 12158 10548 12164 10600
rect 12216 10588 12222 10600
rect 12986 10588 12992 10600
rect 12216 10560 12992 10588
rect 12216 10548 12222 10560
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 13504 10560 17509 10588
rect 13504 10548 13510 10560
rect 17497 10557 17509 10560
rect 17543 10588 17555 10591
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 17543 10560 18521 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 12618 10520 12624 10532
rect 8588 10492 12624 10520
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 14182 10480 14188 10532
rect 14240 10520 14246 10532
rect 17034 10520 17040 10532
rect 14240 10492 17040 10520
rect 14240 10480 14246 10492
rect 17034 10480 17040 10492
rect 17092 10480 17098 10532
rect 10042 10452 10048 10464
rect 8404 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 10284 10424 11529 10452
rect 10284 10412 10290 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 14642 10452 14648 10464
rect 11756 10424 14648 10452
rect 11756 10412 11762 10424
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 16022 10452 16028 10464
rect 14792 10424 16028 10452
rect 14792 10412 14798 10424
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16206 10412 16212 10464
rect 16264 10452 16270 10464
rect 16393 10455 16451 10461
rect 16393 10452 16405 10455
rect 16264 10424 16405 10452
rect 16264 10412 16270 10424
rect 16393 10421 16405 10424
rect 16439 10421 16451 10455
rect 16393 10415 16451 10421
rect 1104 10362 18860 10384
rect 1104 10310 3169 10362
rect 3221 10310 3233 10362
rect 3285 10310 3297 10362
rect 3349 10310 3361 10362
rect 3413 10310 3425 10362
rect 3477 10310 7608 10362
rect 7660 10310 7672 10362
rect 7724 10310 7736 10362
rect 7788 10310 7800 10362
rect 7852 10310 7864 10362
rect 7916 10310 12047 10362
rect 12099 10310 12111 10362
rect 12163 10310 12175 10362
rect 12227 10310 12239 10362
rect 12291 10310 12303 10362
rect 12355 10310 16486 10362
rect 16538 10310 16550 10362
rect 16602 10310 16614 10362
rect 16666 10310 16678 10362
rect 16730 10310 16742 10362
rect 16794 10310 18860 10362
rect 1104 10288 18860 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 3145 10251 3203 10257
rect 3145 10248 3157 10251
rect 1452 10220 3157 10248
rect 1452 10208 1458 10220
rect 3145 10217 3157 10220
rect 3191 10217 3203 10251
rect 3145 10211 3203 10217
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 4798 10248 4804 10260
rect 3651 10220 4804 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 1946 10140 1952 10192
rect 2004 10140 2010 10192
rect 2130 10140 2136 10192
rect 2188 10180 2194 10192
rect 3620 10180 3648 10211
rect 4798 10208 4804 10220
rect 4856 10248 4862 10260
rect 5442 10248 5448 10260
rect 4856 10220 5448 10248
rect 4856 10208 4862 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5902 10248 5908 10260
rect 5592 10220 5908 10248
rect 5592 10208 5598 10220
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 6638 10248 6644 10260
rect 6319 10220 6644 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 2188 10152 3648 10180
rect 2188 10140 2194 10152
rect 3694 10140 3700 10192
rect 3752 10180 3758 10192
rect 4617 10183 4675 10189
rect 4617 10180 4629 10183
rect 3752 10152 4629 10180
rect 3752 10140 3758 10152
rect 4617 10149 4629 10152
rect 4663 10149 4675 10183
rect 4617 10143 4675 10149
rect 4709 10183 4767 10189
rect 4709 10149 4721 10183
rect 4755 10149 4767 10183
rect 6288 10180 6316 10211
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 8202 10248 8208 10260
rect 7800 10220 8208 10248
rect 7800 10208 7806 10220
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 8628 10220 8984 10248
rect 8628 10208 8634 10220
rect 4709 10143 4767 10149
rect 5920 10152 6316 10180
rect 1854 10112 1860 10124
rect 1596 10084 1860 10112
rect 1596 10053 1624 10084
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 1964 10112 1992 10140
rect 1964 10084 2176 10112
rect 2148 10056 2176 10084
rect 2958 10072 2964 10124
rect 3016 10112 3022 10124
rect 4724 10112 4752 10143
rect 5920 10121 5948 10152
rect 7190 10140 7196 10192
rect 7248 10180 7254 10192
rect 8846 10180 8852 10192
rect 7248 10152 8852 10180
rect 7248 10140 7254 10152
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 8956 10180 8984 10220
rect 9306 10208 9312 10260
rect 9364 10208 9370 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 11974 10248 11980 10260
rect 9732 10220 11980 10248
rect 9732 10208 9738 10220
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12176 10220 12388 10248
rect 9398 10180 9404 10192
rect 8956 10152 9404 10180
rect 9398 10140 9404 10152
rect 9456 10140 9462 10192
rect 10778 10140 10784 10192
rect 10836 10140 10842 10192
rect 11054 10140 11060 10192
rect 11112 10180 11118 10192
rect 11701 10183 11759 10189
rect 11701 10180 11713 10183
rect 11112 10152 11713 10180
rect 11112 10140 11118 10152
rect 11701 10149 11713 10152
rect 11747 10180 11759 10183
rect 12176 10180 12204 10220
rect 11747 10152 12204 10180
rect 12360 10180 12388 10220
rect 13906 10208 13912 10260
rect 13964 10208 13970 10260
rect 15746 10248 15752 10260
rect 14016 10220 15752 10248
rect 14016 10180 14044 10220
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 16080 10220 17080 10248
rect 16080 10208 16086 10220
rect 12360 10152 14044 10180
rect 11747 10149 11759 10152
rect 11701 10143 11759 10149
rect 3016 10084 4752 10112
rect 4801 10115 4859 10121
rect 3016 10072 3022 10084
rect 4801 10081 4813 10115
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 1946 10004 1952 10056
rect 2004 10004 2010 10056
rect 2130 10004 2136 10056
rect 2188 10004 2194 10056
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 4154 10044 4160 10056
rect 2915 10016 4160 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 4522 10044 4528 10056
rect 4295 10016 4528 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9976 1915 9979
rect 2406 9976 2412 9988
rect 1903 9948 2412 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 2406 9936 2412 9948
rect 2464 9936 2470 9988
rect 2593 9979 2651 9985
rect 2593 9945 2605 9979
rect 2639 9976 2651 9979
rect 2682 9976 2688 9988
rect 2639 9948 2688 9976
rect 2639 9945 2651 9948
rect 2593 9939 2651 9945
rect 2682 9936 2688 9948
rect 2740 9936 2746 9988
rect 3050 9936 3056 9988
rect 3108 9976 3114 9988
rect 4816 9976 4844 10075
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 6546 10112 6552 10124
rect 6328 10084 6552 10112
rect 6328 10072 6334 10084
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 12158 10112 12164 10124
rect 7340 10084 9674 10112
rect 7340 10072 7346 10084
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 6178 10044 6184 10056
rect 5592 10016 6184 10044
rect 5592 10004 5598 10016
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 7374 10004 7380 10056
rect 7432 10044 7438 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 7432 10016 7481 10044
rect 7432 10004 7438 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7665 10047 7723 10053
rect 7665 10013 7677 10047
rect 7711 10044 7723 10047
rect 8202 10044 8208 10056
rect 7711 10016 8208 10044
rect 7711 10013 7723 10016
rect 7665 10007 7723 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 9364 10016 9505 10044
rect 9364 10004 9370 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9646 10044 9674 10084
rect 10980 10084 12164 10112
rect 10980 10044 11008 10084
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 14826 10112 14832 10124
rect 12268 10084 14832 10112
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 9646 10016 11008 10044
rect 11072 10016 11345 10044
rect 9493 10007 9551 10013
rect 3108 9948 4844 9976
rect 3108 9936 3114 9948
rect 4982 9936 4988 9988
rect 5040 9976 5046 9988
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 5040 9948 5641 9976
rect 5040 9936 5046 9948
rect 5629 9945 5641 9948
rect 5675 9976 5687 9979
rect 8297 9979 8355 9985
rect 8297 9976 8309 9979
rect 5675 9948 8309 9976
rect 5675 9945 5687 9948
rect 5629 9939 5687 9945
rect 8297 9945 8309 9948
rect 8343 9976 8355 9979
rect 9674 9976 9680 9988
rect 8343 9948 9680 9976
rect 8343 9945 8355 9948
rect 8297 9939 8355 9945
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 10962 9936 10968 9988
rect 11020 9976 11026 9988
rect 11072 9976 11100 10016
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11664 10016 11713 10044
rect 11664 10004 11670 10016
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12268 10044 12296 10084
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 14918 10072 14924 10124
rect 14976 10072 14982 10124
rect 12032 10016 12296 10044
rect 12437 10047 12495 10053
rect 12032 10004 12038 10016
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 13170 10044 13176 10056
rect 12667 10016 13176 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 12452 9976 12480 10007
rect 13170 10004 13176 10016
rect 13228 10044 13234 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 13228 10016 13277 10044
rect 13228 10004 13234 10016
rect 13265 10013 13277 10016
rect 13311 10044 13323 10047
rect 14642 10044 14648 10056
rect 13311 10016 14648 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 14936 10044 14964 10072
rect 14936 10016 15042 10044
rect 16390 10004 16396 10056
rect 16448 10004 16454 10056
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 17052 10044 17080 10220
rect 17221 10115 17279 10121
rect 17221 10081 17233 10115
rect 17267 10112 17279 10115
rect 19426 10112 19432 10124
rect 17267 10084 19432 10112
rect 17267 10081 17279 10084
rect 17221 10075 17279 10081
rect 19426 10072 19432 10084
rect 19484 10072 19490 10124
rect 17313 10047 17371 10053
rect 17313 10044 17325 10047
rect 17052 10016 17325 10044
rect 16945 10007 17003 10013
rect 17313 10013 17325 10016
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 12897 9979 12955 9985
rect 12897 9976 12909 9979
rect 11020 9948 11100 9976
rect 12176 9948 12909 9976
rect 11020 9936 11026 9948
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 3786 9908 3792 9920
rect 3660 9880 3792 9908
rect 3660 9868 3666 9880
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 3970 9868 3976 9920
rect 4028 9908 4034 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 4028 9880 4077 9908
rect 4028 9868 4034 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 5077 9911 5135 9917
rect 5077 9908 5089 9911
rect 4764 9880 5089 9908
rect 4764 9868 4770 9880
rect 5077 9877 5089 9880
rect 5123 9877 5135 9911
rect 5077 9871 5135 9877
rect 5353 9911 5411 9917
rect 5353 9877 5365 9911
rect 5399 9908 5411 9911
rect 5442 9908 5448 9920
rect 5399 9880 5448 9908
rect 5399 9877 5411 9880
rect 5353 9871 5411 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 5534 9868 5540 9920
rect 5592 9868 5598 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 5776 9880 6653 9908
rect 5776 9868 5782 9880
rect 6641 9877 6653 9880
rect 6687 9908 6699 9911
rect 9582 9908 9588 9920
rect 6687 9880 9588 9908
rect 6687 9877 6699 9880
rect 6641 9871 6699 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 11238 9908 11244 9920
rect 10928 9880 11244 9908
rect 10928 9868 10934 9880
rect 11238 9868 11244 9880
rect 11296 9908 11302 9920
rect 12176 9908 12204 9948
rect 12897 9945 12909 9948
rect 12943 9976 12955 9979
rect 13446 9976 13452 9988
rect 12943 9948 13452 9976
rect 12943 9945 12955 9948
rect 12897 9939 12955 9945
rect 13446 9936 13452 9948
rect 13504 9936 13510 9988
rect 14369 9979 14427 9985
rect 14369 9945 14381 9979
rect 14415 9976 14427 9979
rect 14458 9976 14464 9988
rect 14415 9948 14464 9976
rect 14415 9945 14427 9948
rect 14369 9939 14427 9945
rect 14458 9936 14464 9948
rect 14516 9936 14522 9988
rect 16117 9979 16175 9985
rect 16117 9945 16129 9979
rect 16163 9976 16175 9979
rect 16850 9976 16856 9988
rect 16163 9948 16856 9976
rect 16163 9945 16175 9948
rect 16117 9939 16175 9945
rect 16850 9936 16856 9948
rect 16908 9936 16914 9988
rect 11296 9880 12204 9908
rect 12253 9911 12311 9917
rect 11296 9868 11302 9880
rect 12253 9877 12265 9911
rect 12299 9908 12311 9911
rect 12342 9908 12348 9920
rect 12299 9880 12348 9908
rect 12299 9877 12311 9880
rect 12253 9871 12311 9877
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 13262 9868 13268 9920
rect 13320 9908 13326 9920
rect 16206 9908 16212 9920
rect 13320 9880 16212 9908
rect 13320 9868 13326 9880
rect 16206 9868 16212 9880
rect 16264 9908 16270 9920
rect 16960 9908 16988 10007
rect 17402 10004 17408 10056
rect 17460 10044 17466 10056
rect 17589 10047 17647 10053
rect 17589 10044 17601 10047
rect 17460 10016 17601 10044
rect 17460 10004 17466 10016
rect 17589 10013 17601 10016
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 17954 10004 17960 10056
rect 18012 10004 18018 10056
rect 16264 9880 16988 9908
rect 16264 9868 16270 9880
rect 1104 9818 18860 9840
rect 1104 9766 3829 9818
rect 3881 9766 3893 9818
rect 3945 9766 3957 9818
rect 4009 9766 4021 9818
rect 4073 9766 4085 9818
rect 4137 9766 8268 9818
rect 8320 9766 8332 9818
rect 8384 9766 8396 9818
rect 8448 9766 8460 9818
rect 8512 9766 8524 9818
rect 8576 9766 12707 9818
rect 12759 9766 12771 9818
rect 12823 9766 12835 9818
rect 12887 9766 12899 9818
rect 12951 9766 12963 9818
rect 13015 9766 17146 9818
rect 17198 9766 17210 9818
rect 17262 9766 17274 9818
rect 17326 9766 17338 9818
rect 17390 9766 17402 9818
rect 17454 9766 18860 9818
rect 1104 9744 18860 9766
rect 2038 9664 2044 9716
rect 2096 9704 2102 9716
rect 2096 9676 3004 9704
rect 2096 9664 2102 9676
rect 1673 9639 1731 9645
rect 1673 9605 1685 9639
rect 1719 9636 1731 9639
rect 1762 9636 1768 9648
rect 1719 9608 1768 9636
rect 1719 9605 1731 9608
rect 1673 9599 1731 9605
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 2682 9596 2688 9648
rect 2740 9596 2746 9648
rect 2976 9636 3004 9676
rect 3602 9664 3608 9716
rect 3660 9704 3666 9716
rect 3786 9704 3792 9716
rect 3660 9676 3792 9704
rect 3660 9664 3666 9676
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7466 9704 7472 9716
rect 7156 9676 7472 9704
rect 7156 9664 7162 9676
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 8941 9707 8999 9713
rect 7576 9676 8892 9704
rect 7576 9648 7604 9676
rect 3697 9639 3755 9645
rect 3697 9636 3709 9639
rect 2976 9608 3709 9636
rect 3697 9605 3709 9608
rect 3743 9605 3755 9639
rect 3697 9599 3755 9605
rect 4801 9639 4859 9645
rect 4801 9605 4813 9639
rect 4847 9636 4859 9639
rect 5626 9636 5632 9648
rect 4847 9608 5632 9636
rect 4847 9605 4859 9608
rect 4801 9599 4859 9605
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 7558 9636 7564 9648
rect 6604 9608 7564 9636
rect 6604 9596 6610 9608
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 8202 9596 8208 9648
rect 8260 9596 8266 9648
rect 8864 9636 8892 9676
rect 8941 9673 8953 9707
rect 8987 9704 8999 9707
rect 9398 9704 9404 9716
rect 8987 9676 9404 9704
rect 8987 9673 8999 9676
rect 8941 9667 8999 9673
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 10226 9704 10232 9716
rect 9732 9676 10232 9704
rect 9732 9664 9738 9676
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 10686 9674 10692 9716
rect 10612 9664 10692 9674
rect 10744 9664 10750 9716
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 13262 9704 13268 9716
rect 11020 9676 13268 9704
rect 11020 9664 11026 9676
rect 10502 9636 10508 9648
rect 8864 9608 10508 9636
rect 10502 9596 10508 9608
rect 10560 9596 10566 9648
rect 10612 9646 10732 9664
rect 3418 9528 3424 9580
rect 3476 9528 3482 9580
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4120 9540 4660 9568
rect 4120 9528 4126 9540
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 1412 9364 1440 9463
rect 4522 9460 4528 9512
rect 4580 9460 4586 9512
rect 4632 9500 4660 9540
rect 4982 9528 4988 9580
rect 5040 9568 5046 9580
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 5040 9540 5089 9568
rect 5040 9528 5046 9540
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 7098 9568 7104 9580
rect 6236 9540 7104 9568
rect 6236 9528 6242 9540
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9674 9568 9680 9580
rect 9364 9540 9680 9568
rect 9364 9528 9370 9540
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 10612 9568 10640 9646
rect 11072 9577 11100 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 13817 9707 13875 9713
rect 11238 9636 11244 9648
rect 11164 9608 11244 9636
rect 11164 9577 11192 9608
rect 11238 9596 11244 9608
rect 11296 9636 11302 9648
rect 11517 9639 11575 9645
rect 11296 9608 11468 9636
rect 11296 9596 11302 9608
rect 10764 9571 10822 9577
rect 10764 9568 10776 9571
rect 10612 9540 10776 9568
rect 10764 9537 10776 9540
rect 10810 9537 10822 9571
rect 10764 9531 10822 9537
rect 10913 9571 10971 9577
rect 10913 9537 10925 9571
rect 10959 9537 10971 9571
rect 10913 9531 10971 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 6638 9500 6644 9512
rect 4632 9472 6644 9500
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 7190 9460 7196 9512
rect 7248 9460 7254 9512
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 8662 9500 8668 9512
rect 7515 9472 8668 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 8846 9460 8852 9512
rect 8904 9500 8910 9512
rect 10226 9500 10232 9512
rect 8904 9472 10232 9500
rect 8904 9460 8910 9472
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 10928 9500 10956 9531
rect 10560 9472 10956 9500
rect 10560 9460 10566 9472
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 4540 9432 4568 9460
rect 4982 9432 4988 9444
rect 4203 9404 4988 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 4982 9392 4988 9404
rect 5040 9392 5046 9444
rect 9493 9435 9551 9441
rect 9493 9401 9505 9435
rect 9539 9432 9551 9435
rect 9674 9432 9680 9444
rect 9539 9404 9680 9432
rect 9539 9401 9551 9404
rect 9493 9395 9551 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9432 9919 9435
rect 11348 9432 11376 9531
rect 11440 9500 11468 9608
rect 11517 9605 11529 9639
rect 11563 9636 11575 9639
rect 11790 9636 11796 9648
rect 11563 9608 11796 9636
rect 11563 9605 11575 9608
rect 11517 9599 11575 9605
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13556 9646 13768 9674
rect 13817 9673 13829 9707
rect 13863 9704 13875 9707
rect 13863 9676 13952 9704
rect 13863 9673 13875 9676
rect 13817 9667 13875 9673
rect 13556 9636 13584 9646
rect 13044 9608 13584 9636
rect 13044 9596 13050 9608
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 11664 9540 12190 9568
rect 13630 9552 13636 9604
rect 13688 9552 13694 9604
rect 11664 9528 11670 9540
rect 13633 9537 13645 9552
rect 13679 9537 13691 9552
rect 13633 9531 13691 9537
rect 13262 9500 13268 9512
rect 11440 9472 13268 9500
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 13538 9460 13544 9512
rect 13596 9460 13602 9512
rect 9907 9404 11376 9432
rect 13740 9432 13768 9646
rect 13924 9580 13952 9676
rect 14090 9664 14096 9716
rect 14148 9664 14154 9716
rect 14366 9664 14372 9716
rect 14424 9704 14430 9716
rect 14424 9676 14872 9704
rect 14424 9664 14430 9676
rect 14292 9608 14688 9636
rect 13906 9528 13912 9580
rect 13964 9528 13970 9580
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14292 9577 14320 9608
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 14056 9540 14289 9568
rect 14056 9528 14062 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14553 9571 14611 9577
rect 14553 9537 14565 9571
rect 14599 9537 14611 9571
rect 14553 9531 14611 9537
rect 14090 9460 14096 9512
rect 14148 9460 14154 9512
rect 14568 9432 14596 9531
rect 13740 9404 14596 9432
rect 14660 9432 14688 9608
rect 14844 9568 14872 9676
rect 16022 9664 16028 9716
rect 16080 9704 16086 9716
rect 16206 9704 16212 9716
rect 16080 9676 16212 9704
rect 16080 9664 16086 9676
rect 16206 9664 16212 9676
rect 16264 9704 16270 9716
rect 17954 9704 17960 9716
rect 16264 9676 17960 9704
rect 16264 9664 16270 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 16298 9596 16304 9648
rect 16356 9636 16362 9648
rect 16356 9608 17724 9636
rect 16356 9596 16362 9608
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14844 9540 14933 9568
rect 14921 9537 14933 9540
rect 14967 9537 14979 9571
rect 16725 9571 16783 9577
rect 16725 9568 16737 9571
rect 14921 9531 14979 9537
rect 16316 9540 16737 9568
rect 16316 9512 16344 9540
rect 16725 9537 16737 9540
rect 16771 9537 16783 9571
rect 16725 9531 16783 9537
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 17696 9577 17724 9608
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 17000 9540 17141 9568
rect 17000 9528 17006 9540
rect 17129 9537 17141 9540
rect 17175 9568 17187 9571
rect 17681 9571 17739 9577
rect 17175 9540 17632 9568
rect 17175 9537 17187 9540
rect 17129 9531 17187 9537
rect 15105 9503 15163 9509
rect 15105 9469 15117 9503
rect 15151 9500 15163 9503
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15151 9472 15393 9500
rect 15151 9469 15163 9472
rect 15105 9463 15163 9469
rect 15381 9469 15393 9472
rect 15427 9500 15439 9503
rect 15654 9500 15660 9512
rect 15427 9472 15660 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 16298 9460 16304 9512
rect 16356 9460 16362 9512
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 16829 9503 16887 9509
rect 16829 9500 16841 9503
rect 16540 9472 16841 9500
rect 16540 9460 16546 9472
rect 16829 9469 16841 9472
rect 16875 9469 16887 9503
rect 16829 9463 16887 9469
rect 17310 9460 17316 9512
rect 17368 9460 17374 9512
rect 15749 9435 15807 9441
rect 15749 9432 15761 9435
rect 14660 9404 15761 9432
rect 9907 9401 9919 9404
rect 9861 9395 9919 9401
rect 15749 9401 15761 9404
rect 15795 9432 15807 9435
rect 15930 9432 15936 9444
rect 15795 9404 15936 9432
rect 15795 9401 15807 9404
rect 15749 9395 15807 9401
rect 3510 9364 3516 9376
rect 1412 9336 3516 9364
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 4580 9336 5549 9364
rect 4580 9324 4586 9336
rect 5537 9333 5549 9336
rect 5583 9364 5595 9367
rect 6638 9364 6644 9376
rect 5583 9336 6644 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 8202 9364 8208 9376
rect 7156 9336 8208 9364
rect 7156 9324 7162 9336
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 9582 9324 9588 9376
rect 9640 9364 9646 9376
rect 9876 9364 9904 9395
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 9640 9336 9904 9364
rect 9640 9324 9646 9336
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 10560 9336 10609 9364
rect 10560 9324 10566 9336
rect 10597 9333 10609 9336
rect 10643 9364 10655 9367
rect 11054 9364 11060 9376
rect 10643 9336 11060 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 11974 9364 11980 9376
rect 11848 9336 11980 9364
rect 11848 9324 11854 9336
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13277 9367 13335 9373
rect 13277 9364 13289 9367
rect 13136 9336 13289 9364
rect 13136 9324 13142 9336
rect 13277 9333 13289 9336
rect 13323 9333 13335 9367
rect 13277 9327 13335 9333
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 15378 9364 15384 9376
rect 14424 9336 15384 9364
rect 14424 9324 14430 9336
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 16206 9324 16212 9376
rect 16264 9324 16270 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17034 9364 17040 9376
rect 16816 9336 17040 9364
rect 16816 9324 16822 9336
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 17126 9324 17132 9376
rect 17184 9364 17190 9376
rect 17497 9367 17555 9373
rect 17497 9364 17509 9367
rect 17184 9336 17509 9364
rect 17184 9324 17190 9336
rect 17497 9333 17509 9336
rect 17543 9333 17555 9367
rect 17604 9364 17632 9540
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 17773 9571 17831 9577
rect 17773 9537 17785 9571
rect 17819 9568 17831 9571
rect 18414 9568 18420 9580
rect 17819 9540 18420 9568
rect 17819 9537 17831 9540
rect 17773 9531 17831 9537
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17920 9472 18061 9500
rect 17920 9460 17926 9472
rect 18049 9469 18061 9472
rect 18095 9500 18107 9503
rect 18325 9503 18383 9509
rect 18325 9500 18337 9503
rect 18095 9472 18337 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18325 9469 18337 9472
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 17957 9367 18015 9373
rect 17957 9364 17969 9367
rect 17604 9336 17969 9364
rect 17497 9327 17555 9333
rect 17957 9333 17969 9336
rect 18003 9364 18015 9367
rect 18506 9364 18512 9376
rect 18003 9336 18512 9364
rect 18003 9333 18015 9336
rect 17957 9327 18015 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 1104 9274 18860 9296
rect 1104 9222 3169 9274
rect 3221 9222 3233 9274
rect 3285 9222 3297 9274
rect 3349 9222 3361 9274
rect 3413 9222 3425 9274
rect 3477 9222 7608 9274
rect 7660 9222 7672 9274
rect 7724 9222 7736 9274
rect 7788 9222 7800 9274
rect 7852 9222 7864 9274
rect 7916 9222 12047 9274
rect 12099 9222 12111 9274
rect 12163 9222 12175 9274
rect 12227 9222 12239 9274
rect 12291 9222 12303 9274
rect 12355 9222 16486 9274
rect 16538 9222 16550 9274
rect 16602 9222 16614 9274
rect 16666 9222 16678 9274
rect 16730 9222 16742 9274
rect 16794 9222 18860 9274
rect 1104 9200 18860 9222
rect 2314 9120 2320 9172
rect 2372 9120 2378 9172
rect 2501 9163 2559 9169
rect 2501 9129 2513 9163
rect 2547 9160 2559 9163
rect 2590 9160 2596 9172
rect 2547 9132 2596 9160
rect 2547 9129 2559 9132
rect 2501 9123 2559 9129
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 2866 9120 2872 9172
rect 2924 9120 2930 9172
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4154 9160 4160 9172
rect 3844 9132 4160 9160
rect 3844 9120 3850 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 5261 9163 5319 9169
rect 5261 9160 5273 9163
rect 4396 9132 5273 9160
rect 4396 9120 4402 9132
rect 5261 9129 5273 9132
rect 5307 9160 5319 9163
rect 5442 9160 5448 9172
rect 5307 9132 5448 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 5442 9120 5448 9132
rect 5500 9160 5506 9172
rect 6086 9160 6092 9172
rect 5500 9132 6092 9160
rect 5500 9120 5506 9132
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 6181 9163 6239 9169
rect 6181 9129 6193 9163
rect 6227 9160 6239 9163
rect 6914 9160 6920 9172
rect 6227 9132 6920 9160
rect 6227 9129 6239 9132
rect 6181 9123 6239 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 7800 9132 8708 9160
rect 7800 9120 7806 9132
rect 2222 9052 2228 9104
rect 2280 9052 2286 9104
rect 3602 9052 3608 9104
rect 3660 9092 3666 9104
rect 7006 9092 7012 9104
rect 3660 9064 7012 9092
rect 3660 9052 3666 9064
rect 7006 9052 7012 9064
rect 7064 9052 7070 9104
rect 8680 9092 8708 9132
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 10318 9160 10324 9172
rect 9732 9132 10324 9160
rect 9732 9120 9738 9132
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 10686 9120 10692 9172
rect 10744 9160 10750 9172
rect 13814 9160 13820 9172
rect 10744 9132 13820 9160
rect 10744 9120 10750 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 15197 9163 15255 9169
rect 15197 9160 15209 9163
rect 14884 9132 15209 9160
rect 14884 9120 14890 9132
rect 15197 9129 15209 9132
rect 15243 9160 15255 9163
rect 15378 9160 15384 9172
rect 15243 9132 15384 9160
rect 15243 9129 15255 9132
rect 15197 9123 15255 9129
rect 15378 9120 15384 9132
rect 15436 9160 15442 9172
rect 15654 9160 15660 9172
rect 15436 9132 15660 9160
rect 15436 9120 15442 9132
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 15749 9163 15807 9169
rect 15749 9129 15761 9163
rect 15795 9160 15807 9163
rect 16022 9160 16028 9172
rect 15795 9132 16028 9160
rect 15795 9129 15807 9132
rect 15749 9123 15807 9129
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 17310 9160 17316 9172
rect 16316 9132 17316 9160
rect 10962 9092 10968 9104
rect 8680 9064 10968 9092
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 11149 9095 11207 9101
rect 11149 9092 11161 9095
rect 11072 9064 11161 9092
rect 2240 9024 2268 9052
rect 2240 8996 2774 9024
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2409 8959 2467 8965
rect 2409 8956 2421 8959
rect 2280 8928 2421 8956
rect 2280 8916 2286 8928
rect 2409 8925 2421 8928
rect 2455 8925 2467 8959
rect 2746 8956 2774 8996
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 2924 8996 4629 9024
rect 2924 8984 2930 8996
rect 4617 8993 4629 8996
rect 4663 9024 4675 9027
rect 5626 9024 5632 9036
rect 4663 8996 5632 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5767 8996 5825 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 5813 8993 5825 8996
rect 5859 9024 5871 9027
rect 6914 9024 6920 9036
rect 5859 8996 6920 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 8386 9024 8392 9036
rect 7892 8996 8392 9024
rect 7892 8984 7898 8996
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 10686 9024 10692 9036
rect 8527 8996 10692 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 3234 8956 3240 8968
rect 2746 8928 3240 8956
rect 2409 8919 2467 8925
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 4430 8956 4436 8968
rect 4387 8928 4436 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5500 8928 6009 8956
rect 5500 8916 5506 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 7098 8956 7104 8968
rect 5997 8919 6055 8925
rect 6104 8928 7104 8956
rect 2038 8848 2044 8900
rect 2096 8888 2102 8900
rect 2096 8860 4844 8888
rect 2096 8848 2102 8860
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3973 8823 4031 8829
rect 3973 8820 3985 8823
rect 3108 8792 3985 8820
rect 3108 8780 3114 8792
rect 3973 8789 3985 8792
rect 4019 8789 4031 8823
rect 3973 8783 4031 8789
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 4522 8820 4528 8832
rect 4479 8792 4528 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4816 8820 4844 8860
rect 5626 8848 5632 8900
rect 5684 8888 5690 8900
rect 6104 8888 6132 8928
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 8754 8916 8760 8968
rect 8812 8916 8818 8968
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9582 8916 9588 8968
rect 9640 8916 9646 8968
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9824 8928 9965 8956
rect 9824 8916 9830 8928
rect 9953 8925 9965 8928
rect 9999 8956 10011 8959
rect 10134 8956 10140 8968
rect 9999 8928 10140 8956
rect 9999 8925 10011 8928
rect 9953 8919 10011 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10318 8916 10324 8968
rect 10376 8916 10382 8968
rect 11072 8956 11100 9064
rect 11149 9061 11161 9064
rect 11195 9092 11207 9095
rect 11514 9092 11520 9104
rect 11195 9064 11520 9092
rect 11195 9061 11207 9064
rect 11149 9055 11207 9061
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 16316 9092 16344 9132
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 12924 9064 13768 9092
rect 12924 9024 12952 9064
rect 10428 8928 11100 8956
rect 11440 8996 12952 9024
rect 5684 8860 6132 8888
rect 6273 8891 6331 8897
rect 5684 8848 5690 8860
rect 6273 8857 6285 8891
rect 6319 8888 6331 8891
rect 7190 8888 7196 8900
rect 6319 8860 7196 8888
rect 6319 8857 6331 8860
rect 6273 8851 6331 8857
rect 7190 8848 7196 8860
rect 7248 8848 7254 8900
rect 8202 8888 8208 8900
rect 8050 8860 8208 8888
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 9232 8888 9260 8916
rect 10428 8888 10456 8928
rect 9232 8860 10456 8888
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 4816 8792 7021 8820
rect 7009 8789 7021 8792
rect 7055 8820 7067 8823
rect 11440 8820 11468 8996
rect 12986 8984 12992 9036
rect 13044 8984 13050 9036
rect 13357 9027 13415 9033
rect 13357 8993 13369 9027
rect 13403 9024 13415 9027
rect 13538 9024 13544 9036
rect 13403 8996 13544 9024
rect 13403 8993 13415 8996
rect 13357 8987 13415 8993
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 13740 9024 13768 9064
rect 16040 9064 16344 9092
rect 16040 9033 16068 9064
rect 16390 9052 16396 9104
rect 16448 9052 16454 9104
rect 16025 9027 16083 9033
rect 16025 9024 16037 9027
rect 13740 8996 16037 9024
rect 16025 8993 16037 8996
rect 16071 8993 16083 9027
rect 16408 9024 16436 9052
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16408 8996 16497 9024
rect 16025 8987 16083 8993
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 16758 8984 16764 9036
rect 16816 9024 16822 9036
rect 17954 9024 17960 9036
rect 16816 8996 17960 9024
rect 16816 8984 16822 8996
rect 17954 8984 17960 8996
rect 18012 9024 18018 9036
rect 18233 9027 18291 9033
rect 18233 9024 18245 9027
rect 18012 8996 18245 9024
rect 18012 8984 18018 8996
rect 18233 8993 18245 8996
rect 18279 8993 18291 9027
rect 18233 8987 18291 8993
rect 11606 8916 11612 8968
rect 11664 8956 11670 8968
rect 12529 8959 12587 8965
rect 11664 8928 11836 8956
rect 11664 8916 11670 8928
rect 11808 8900 11836 8928
rect 12529 8925 12541 8959
rect 12575 8956 12587 8959
rect 12618 8956 12624 8968
rect 12575 8928 12624 8956
rect 12575 8925 12587 8928
rect 12529 8919 12587 8925
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8956 12955 8959
rect 13630 8956 13636 8968
rect 12943 8928 13636 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13872 8928 14105 8956
rect 13872 8916 13878 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 15010 8916 15016 8968
rect 15068 8956 15074 8968
rect 16298 8956 16304 8968
rect 15068 8928 16304 8956
rect 15068 8916 15074 8928
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16390 8916 16396 8968
rect 16448 8916 16454 8968
rect 11790 8848 11796 8900
rect 11848 8848 11854 8900
rect 13449 8891 13507 8897
rect 13449 8857 13461 8891
rect 13495 8857 13507 8891
rect 13449 8851 13507 8857
rect 13725 8891 13783 8897
rect 13725 8857 13737 8891
rect 13771 8888 13783 8891
rect 15102 8888 15108 8900
rect 13771 8860 15108 8888
rect 13771 8857 13783 8860
rect 13725 8851 13783 8857
rect 7055 8792 11468 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 11606 8780 11612 8832
rect 11664 8820 11670 8832
rect 12618 8820 12624 8832
rect 11664 8792 12624 8820
rect 11664 8780 11670 8792
rect 12618 8780 12624 8792
rect 12676 8820 12682 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 12676 8792 13277 8820
rect 12676 8780 12682 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13469 8820 13497 8851
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 16022 8888 16028 8900
rect 15528 8860 16028 8888
rect 15528 8848 15534 8860
rect 16022 8848 16028 8860
rect 16080 8848 16086 8900
rect 16761 8891 16819 8897
rect 16761 8857 16773 8891
rect 16807 8857 16819 8891
rect 16761 8851 16819 8857
rect 14182 8820 14188 8832
rect 13469 8792 14188 8820
rect 13265 8783 13323 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14274 8780 14280 8832
rect 14332 8780 14338 8832
rect 14645 8823 14703 8829
rect 14645 8789 14657 8823
rect 14691 8820 14703 8823
rect 14918 8820 14924 8832
rect 14691 8792 14924 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 16209 8823 16267 8829
rect 16209 8789 16221 8823
rect 16255 8820 16267 8823
rect 16298 8820 16304 8832
rect 16255 8792 16304 8820
rect 16255 8789 16267 8792
rect 16209 8783 16267 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 16776 8820 16804 8851
rect 17034 8848 17040 8900
rect 17092 8888 17098 8900
rect 17092 8860 17250 8888
rect 17092 8848 17098 8860
rect 17402 8820 17408 8832
rect 16776 8792 17408 8820
rect 17402 8780 17408 8792
rect 17460 8780 17466 8832
rect 1104 8730 18860 8752
rect 1104 8678 3829 8730
rect 3881 8678 3893 8730
rect 3945 8678 3957 8730
rect 4009 8678 4021 8730
rect 4073 8678 4085 8730
rect 4137 8678 8268 8730
rect 8320 8678 8332 8730
rect 8384 8678 8396 8730
rect 8448 8678 8460 8730
rect 8512 8678 8524 8730
rect 8576 8678 12707 8730
rect 12759 8678 12771 8730
rect 12823 8678 12835 8730
rect 12887 8678 12899 8730
rect 12951 8678 12963 8730
rect 13015 8678 17146 8730
rect 17198 8678 17210 8730
rect 17262 8678 17274 8730
rect 17326 8678 17338 8730
rect 17390 8678 17402 8730
rect 17454 8678 18860 8730
rect 1104 8656 18860 8678
rect 2958 8616 2964 8628
rect 1596 8588 2964 8616
rect 1596 8489 1624 8588
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 3510 8576 3516 8628
rect 3568 8616 3574 8628
rect 3568 8588 5948 8616
rect 3568 8576 3574 8588
rect 3142 8548 3148 8560
rect 1688 8520 3148 8548
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 1688 8421 1716 8520
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 3602 8508 3608 8560
rect 3660 8548 3666 8560
rect 3789 8551 3847 8557
rect 3789 8548 3801 8551
rect 3660 8520 3801 8548
rect 3660 8508 3666 8520
rect 3789 8517 3801 8520
rect 3835 8517 3847 8551
rect 5626 8548 5632 8560
rect 5106 8520 5632 8548
rect 3789 8511 3847 8517
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 3694 8480 3700 8492
rect 2179 8452 3700 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5920 8480 5948 8588
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 8386 8616 8392 8628
rect 6052 8588 8392 8616
rect 6052 8576 6058 8588
rect 8386 8576 8392 8588
rect 8444 8616 8450 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 8444 8588 8953 8616
rect 8444 8576 8450 8588
rect 8941 8585 8953 8588
rect 8987 8616 8999 8619
rect 9490 8616 9496 8628
rect 8987 8588 9496 8616
rect 8987 8585 8999 8588
rect 8941 8579 8999 8585
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 10410 8616 10416 8628
rect 9640 8588 10416 8616
rect 9640 8576 9646 8588
rect 10410 8576 10416 8588
rect 10468 8616 10474 8628
rect 11606 8616 11612 8628
rect 10468 8588 11612 8616
rect 10468 8576 10474 8588
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 13725 8619 13783 8625
rect 13725 8616 13737 8619
rect 12492 8588 13737 8616
rect 12492 8576 12498 8588
rect 13725 8585 13737 8588
rect 13771 8585 13783 8619
rect 13725 8579 13783 8585
rect 13998 8576 14004 8628
rect 14056 8576 14062 8628
rect 15105 8619 15163 8625
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 15838 8616 15844 8628
rect 15151 8588 15844 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 16850 8576 16856 8628
rect 16908 8576 16914 8628
rect 16942 8576 16948 8628
rect 17000 8616 17006 8628
rect 17126 8616 17132 8628
rect 17000 8588 17132 8616
rect 17000 8576 17006 8588
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17218 8576 17224 8628
rect 17276 8616 17282 8628
rect 17678 8616 17684 8628
rect 17276 8588 17684 8616
rect 17276 8576 17282 8588
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 18414 8576 18420 8628
rect 18472 8576 18478 8628
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 7558 8548 7564 8560
rect 7064 8520 7564 8548
rect 7064 8508 7070 8520
rect 7558 8508 7564 8520
rect 7616 8508 7622 8560
rect 8110 8508 8116 8560
rect 8168 8508 8174 8560
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 8846 8548 8852 8560
rect 8536 8520 8852 8548
rect 8536 8508 8542 8520
rect 8846 8508 8852 8520
rect 8904 8508 8910 8560
rect 11146 8508 11152 8560
rect 11204 8548 11210 8560
rect 11517 8551 11575 8557
rect 11517 8548 11529 8551
rect 11204 8520 11529 8548
rect 11204 8508 11210 8520
rect 11517 8517 11529 8520
rect 11563 8517 11575 8551
rect 11517 8511 11575 8517
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 11848 8534 12006 8548
rect 11848 8520 12020 8534
rect 11848 8508 11854 8520
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5859 8452 6377 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6365 8449 6377 8452
rect 6411 8480 6423 8483
rect 7190 8480 7196 8492
rect 6411 8452 7196 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 9306 8480 9312 8492
rect 8812 8452 9312 8480
rect 8812 8440 8818 8452
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8381 1823 8415
rect 1765 8375 1823 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 8662 8412 8668 8424
rect 5583 8384 8668 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 1210 8304 1216 8356
rect 1268 8344 1274 8356
rect 1780 8344 1808 8375
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 8904 8384 9597 8412
rect 8904 8372 8910 8384
rect 9585 8381 9597 8384
rect 9631 8381 9643 8415
rect 10704 8412 10732 8440
rect 11992 8412 12020 8520
rect 15378 8508 15384 8560
rect 15436 8548 15442 8560
rect 15749 8551 15807 8557
rect 15749 8548 15761 8551
rect 15436 8520 15761 8548
rect 15436 8508 15442 8520
rect 15749 8517 15761 8520
rect 15795 8517 15807 8551
rect 18141 8551 18199 8557
rect 18141 8548 18153 8551
rect 15749 8511 15807 8517
rect 15856 8520 17448 8548
rect 12894 8440 12900 8492
rect 12952 8480 12958 8492
rect 15856 8480 15884 8520
rect 16758 8480 16764 8492
rect 12952 8452 15884 8480
rect 15948 8452 16764 8480
rect 12952 8440 12958 8452
rect 12526 8412 12532 8424
rect 10704 8384 12532 8412
rect 9585 8375 9643 8381
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 12676 8384 13001 8412
rect 12676 8372 12682 8384
rect 12989 8381 13001 8384
rect 13035 8381 13047 8415
rect 12989 8375 13047 8381
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8412 13415 8415
rect 13630 8412 13636 8424
rect 13403 8384 13636 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 14182 8372 14188 8424
rect 14240 8412 14246 8424
rect 15948 8412 15976 8452
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17218 8480 17224 8492
rect 17083 8452 17224 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 14240 8384 15976 8412
rect 14240 8372 14246 8384
rect 16022 8372 16028 8424
rect 16080 8372 16086 8424
rect 16390 8412 16396 8424
rect 16132 8384 16396 8412
rect 1268 8316 1808 8344
rect 1268 8304 1274 8316
rect 6086 8304 6092 8356
rect 6144 8344 6150 8356
rect 8478 8344 8484 8356
rect 6144 8316 8484 8344
rect 6144 8304 6150 8316
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 9030 8344 9036 8356
rect 8628 8316 9036 8344
rect 8628 8304 8634 8316
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 11112 8316 12020 8344
rect 11112 8304 11118 8316
rect 11992 8288 12020 8316
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 13596 8316 15240 8344
rect 13596 8304 13602 8316
rect 15212 8288 15240 8316
rect 15378 8304 15384 8356
rect 15436 8304 15442 8356
rect 16132 8344 16160 8384
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 16942 8372 16948 8424
rect 17000 8412 17006 8424
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 17000 8384 17141 8412
rect 17000 8372 17006 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 17310 8372 17316 8424
rect 17368 8372 17374 8424
rect 17420 8344 17448 8520
rect 17696 8520 18153 8548
rect 17696 8492 17724 8520
rect 18141 8517 18153 8520
rect 18187 8517 18199 8551
rect 18141 8511 18199 8517
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 17866 8483 17924 8489
rect 17866 8449 17878 8483
rect 17912 8480 17924 8483
rect 17954 8480 17960 8492
rect 17912 8452 17960 8480
rect 17912 8449 17924 8452
rect 17866 8443 17924 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 18279 8483 18337 8489
rect 18279 8449 18291 8483
rect 18325 8480 18337 8483
rect 18325 8452 18644 8480
rect 18325 8449 18337 8452
rect 18279 8443 18337 8449
rect 17494 8372 17500 8424
rect 17552 8372 17558 8424
rect 18064 8412 18092 8443
rect 18506 8412 18512 8424
rect 18064 8384 18512 8412
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 17770 8344 17776 8356
rect 15488 8316 16160 8344
rect 16316 8316 17172 8344
rect 17420 8316 17776 8344
rect 1854 8236 1860 8288
rect 1912 8276 1918 8288
rect 2409 8279 2467 8285
rect 2409 8276 2421 8279
rect 1912 8248 2421 8276
rect 1912 8236 1918 8248
rect 2409 8245 2421 8248
rect 2455 8245 2467 8279
rect 2409 8239 2467 8245
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3234 8276 3240 8288
rect 3016 8248 3240 8276
rect 3016 8236 3022 8248
rect 3234 8236 3240 8248
rect 3292 8276 3298 8288
rect 3694 8276 3700 8288
rect 3292 8248 3700 8276
rect 3292 8236 3298 8248
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 11330 8276 11336 8288
rect 5040 8248 11336 8276
rect 5040 8236 5046 8248
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 14737 8279 14795 8285
rect 14737 8276 14749 8279
rect 12032 8248 14749 8276
rect 12032 8236 12038 8248
rect 14737 8245 14749 8248
rect 14783 8276 14795 8279
rect 15102 8276 15108 8288
rect 14783 8248 15108 8276
rect 14783 8245 14795 8248
rect 14737 8239 14795 8245
rect 15102 8236 15108 8248
rect 15160 8236 15166 8288
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 15488 8276 15516 8316
rect 15252 8248 15516 8276
rect 15252 8236 15258 8248
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 16316 8276 16344 8316
rect 15896 8248 16344 8276
rect 17144 8276 17172 8316
rect 17770 8304 17776 8316
rect 17828 8344 17834 8356
rect 18616 8344 18644 8452
rect 17828 8316 18644 8344
rect 17828 8304 17834 8316
rect 18966 8276 18972 8288
rect 17144 8248 18972 8276
rect 15896 8236 15902 8248
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 1104 8186 18860 8208
rect 1104 8134 3169 8186
rect 3221 8134 3233 8186
rect 3285 8134 3297 8186
rect 3349 8134 3361 8186
rect 3413 8134 3425 8186
rect 3477 8134 7608 8186
rect 7660 8134 7672 8186
rect 7724 8134 7736 8186
rect 7788 8134 7800 8186
rect 7852 8134 7864 8186
rect 7916 8134 12047 8186
rect 12099 8134 12111 8186
rect 12163 8134 12175 8186
rect 12227 8134 12239 8186
rect 12291 8134 12303 8186
rect 12355 8134 16486 8186
rect 16538 8134 16550 8186
rect 16602 8134 16614 8186
rect 16666 8134 16678 8186
rect 16730 8134 16742 8186
rect 16794 8134 18860 8186
rect 1104 8112 18860 8134
rect 2685 8075 2743 8081
rect 2685 8072 2697 8075
rect 1872 8044 2697 8072
rect 1578 7896 1584 7948
rect 1636 7896 1642 7948
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1762 7868 1768 7880
rect 900 7840 1768 7868
rect 900 7828 906 7840
rect 1762 7828 1768 7840
rect 1820 7868 1826 7880
rect 1872 7877 1900 8044
rect 2685 8041 2697 8044
rect 2731 8041 2743 8075
rect 2685 8035 2743 8041
rect 3145 8075 3203 8081
rect 3145 8041 3157 8075
rect 3191 8072 3203 8075
rect 6178 8072 6184 8084
rect 3191 8044 6184 8072
rect 3191 8041 3203 8044
rect 3145 8035 3203 8041
rect 2130 7964 2136 8016
rect 2188 8004 2194 8016
rect 2590 8004 2596 8016
rect 2188 7976 2596 8004
rect 2188 7964 2194 7976
rect 2590 7964 2596 7976
rect 2648 7964 2654 8016
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 3160 7936 3188 8035
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 6362 8032 6368 8084
rect 6420 8032 6426 8084
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 8570 8072 8576 8084
rect 7156 8044 8576 8072
rect 7156 8032 7162 8044
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 8680 8044 9873 8072
rect 6380 8004 6408 8032
rect 2372 7908 3188 7936
rect 4724 7976 6408 8004
rect 2372 7896 2378 7908
rect 1857 7871 1915 7877
rect 1857 7868 1869 7871
rect 1820 7840 1869 7868
rect 1820 7828 1826 7840
rect 1857 7837 1869 7840
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7868 2467 7871
rect 3602 7868 3608 7880
rect 2455 7840 3608 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 4338 7868 4344 7880
rect 4111 7840 4344 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 4724 7868 4752 7976
rect 8680 7945 8708 8044
rect 9861 8041 9873 8044
rect 9907 8072 9919 8075
rect 12066 8072 12072 8084
rect 9907 8044 12072 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 12526 8072 12532 8084
rect 12308 8044 12532 8072
rect 12308 8032 12314 8044
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13814 8072 13820 8084
rect 13504 8044 13820 8072
rect 13504 8032 13510 8044
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 13909 8075 13967 8081
rect 13909 8041 13921 8075
rect 13955 8072 13967 8075
rect 14366 8072 14372 8084
rect 13955 8044 14372 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 15746 8072 15752 8084
rect 15703 8044 15752 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 16022 8032 16028 8084
rect 16080 8072 16086 8084
rect 16301 8075 16359 8081
rect 16301 8072 16313 8075
rect 16080 8044 16313 8072
rect 16080 8032 16086 8044
rect 16301 8041 16313 8044
rect 16347 8041 16359 8075
rect 16301 8035 16359 8041
rect 16390 8032 16396 8084
rect 16448 8072 16454 8084
rect 17034 8072 17040 8084
rect 16448 8044 17040 8072
rect 16448 8032 16454 8044
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 9125 8007 9183 8013
rect 9125 7973 9137 8007
rect 9171 8004 9183 8007
rect 9171 7976 9674 8004
rect 9171 7973 9183 7976
rect 9125 7967 9183 7973
rect 8665 7939 8723 7945
rect 8665 7936 8677 7939
rect 4908 7908 8677 7936
rect 4479 7840 4752 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 4798 7828 4804 7880
rect 4856 7828 4862 7880
rect 2130 7760 2136 7812
rect 2188 7760 2194 7812
rect 4908 7800 4936 7908
rect 8665 7905 8677 7908
rect 8711 7905 8723 7939
rect 9398 7936 9404 7948
rect 8665 7899 8723 7905
rect 9324 7908 9404 7936
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5132 7840 5549 7868
rect 5132 7828 5138 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 9324 7877 9352 7908
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9490 7896 9496 7948
rect 9548 7896 9554 7948
rect 9646 7936 9674 7976
rect 11330 7964 11336 8016
rect 11388 8004 11394 8016
rect 11388 7976 14964 8004
rect 11388 7964 11394 7976
rect 9858 7936 9864 7948
rect 9646 7908 9864 7936
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 10686 7896 10692 7948
rect 10744 7896 10750 7948
rect 11164 7908 13676 7936
rect 11164 7880 11192 7908
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 8444 7840 9321 7868
rect 8444 7828 8450 7840
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 10965 7871 11023 7877
rect 9309 7831 9367 7837
rect 9600 7840 10916 7868
rect 2240 7772 4936 7800
rect 4985 7803 5043 7809
rect 1302 7692 1308 7744
rect 1360 7732 1366 7744
rect 2240 7732 2268 7772
rect 4985 7769 4997 7803
rect 5031 7800 5043 7803
rect 5442 7800 5448 7812
rect 5031 7772 5448 7800
rect 5031 7769 5043 7772
rect 4985 7763 5043 7769
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 5994 7760 6000 7812
rect 6052 7800 6058 7812
rect 6052 7772 9168 7800
rect 6052 7760 6058 7772
rect 1360 7704 2268 7732
rect 1360 7692 1366 7704
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 5902 7732 5908 7744
rect 4396 7704 5908 7732
rect 4396 7692 4402 7704
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 6822 7692 6828 7744
rect 6880 7732 6886 7744
rect 9030 7732 9036 7744
rect 6880 7704 9036 7732
rect 6880 7692 6886 7704
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9140 7732 9168 7772
rect 9600 7732 9628 7840
rect 10045 7803 10103 7809
rect 10045 7769 10057 7803
rect 10091 7800 10103 7803
rect 10410 7800 10416 7812
rect 10091 7772 10416 7800
rect 10091 7769 10103 7772
rect 10045 7763 10103 7769
rect 10410 7760 10416 7772
rect 10468 7760 10474 7812
rect 10888 7800 10916 7840
rect 10965 7837 10977 7871
rect 11011 7868 11023 7871
rect 11146 7868 11152 7880
rect 11011 7840 11152 7868
rect 11011 7837 11023 7840
rect 10965 7831 11023 7837
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12032 7840 13584 7868
rect 12032 7828 12038 7840
rect 12710 7800 12716 7812
rect 10888 7772 12716 7800
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 9140 7704 9628 7732
rect 9677 7735 9735 7741
rect 9677 7701 9689 7735
rect 9723 7732 9735 7735
rect 9766 7732 9772 7744
rect 9723 7704 9772 7732
rect 9723 7701 9735 7704
rect 9677 7695 9735 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 9861 7735 9919 7741
rect 9861 7701 9873 7735
rect 9907 7732 9919 7735
rect 9950 7732 9956 7744
rect 9907 7704 9956 7732
rect 9907 7701 9919 7704
rect 9861 7695 9919 7701
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 10284 7704 10333 7732
rect 10284 7692 10290 7704
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 10502 7692 10508 7744
rect 10560 7732 10566 7744
rect 10870 7732 10876 7744
rect 10560 7704 10876 7732
rect 10560 7692 10566 7704
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 11330 7692 11336 7744
rect 11388 7732 11394 7744
rect 11514 7732 11520 7744
rect 11388 7704 11520 7732
rect 11388 7692 11394 7704
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 11606 7692 11612 7744
rect 11664 7692 11670 7744
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 12802 7732 12808 7744
rect 12308 7704 12808 7732
rect 12308 7692 12314 7704
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 13556 7732 13584 7840
rect 13648 7800 13676 7908
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 13780 7908 14841 7936
rect 13780 7896 13786 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14936 7936 14964 7976
rect 15010 7964 15016 8016
rect 15068 7964 15074 8016
rect 16761 8007 16819 8013
rect 16761 8004 16773 8007
rect 15120 7976 16773 8004
rect 15120 7936 15148 7976
rect 16761 7973 16773 7976
rect 16807 8004 16819 8007
rect 17310 8004 17316 8016
rect 16807 7976 17316 8004
rect 16807 7973 16819 7976
rect 16761 7967 16819 7973
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 17681 8007 17739 8013
rect 17681 7973 17693 8007
rect 17727 8004 17739 8007
rect 18414 8004 18420 8016
rect 17727 7976 18420 8004
rect 17727 7973 17739 7976
rect 17681 7967 17739 7973
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 14936 7908 15148 7936
rect 14829 7899 14887 7905
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 15620 7908 18276 7936
rect 15620 7896 15626 7908
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 15013 7871 15071 7877
rect 15013 7868 15025 7871
rect 14792 7840 15025 7868
rect 14792 7828 14798 7840
rect 15013 7837 15025 7840
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7868 16083 7871
rect 17313 7871 17371 7877
rect 16071 7840 17264 7868
rect 16071 7837 16083 7840
rect 16025 7831 16083 7837
rect 14918 7800 14924 7812
rect 13648 7772 14924 7800
rect 14918 7760 14924 7772
rect 14976 7760 14982 7812
rect 15102 7760 15108 7812
rect 15160 7800 15166 7812
rect 15381 7803 15439 7809
rect 15381 7800 15393 7803
rect 15160 7772 15393 7800
rect 15160 7760 15166 7772
rect 15381 7769 15393 7772
rect 15427 7800 15439 7803
rect 15562 7800 15568 7812
rect 15427 7772 15568 7800
rect 15427 7769 15439 7772
rect 15381 7763 15439 7769
rect 15562 7760 15568 7772
rect 15620 7760 15626 7812
rect 15672 7800 15700 7831
rect 16850 7800 16856 7812
rect 15672 7772 16856 7800
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 17236 7800 17264 7840
rect 17313 7837 17325 7871
rect 17359 7868 17371 7871
rect 17494 7868 17500 7880
rect 17359 7840 17500 7868
rect 17359 7837 17371 7840
rect 17313 7831 17371 7837
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 18248 7877 18276 7908
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 17236 7772 18276 7800
rect 18248 7744 18276 7772
rect 14090 7732 14096 7744
rect 13556 7704 14096 7732
rect 14090 7692 14096 7704
rect 14148 7732 14154 7744
rect 14277 7735 14335 7741
rect 14277 7732 14289 7735
rect 14148 7704 14289 7732
rect 14148 7692 14154 7704
rect 14277 7701 14289 7704
rect 14323 7701 14335 7735
rect 14277 7695 14335 7701
rect 14734 7692 14740 7744
rect 14792 7692 14798 7744
rect 15838 7692 15844 7744
rect 15896 7692 15902 7744
rect 17126 7692 17132 7744
rect 17184 7692 17190 7744
rect 18046 7692 18052 7744
rect 18104 7692 18110 7744
rect 18230 7692 18236 7744
rect 18288 7692 18294 7744
rect 1104 7642 18860 7664
rect 1104 7590 3829 7642
rect 3881 7590 3893 7642
rect 3945 7590 3957 7642
rect 4009 7590 4021 7642
rect 4073 7590 4085 7642
rect 4137 7590 8268 7642
rect 8320 7590 8332 7642
rect 8384 7590 8396 7642
rect 8448 7590 8460 7642
rect 8512 7590 8524 7642
rect 8576 7590 12707 7642
rect 12759 7590 12771 7642
rect 12823 7590 12835 7642
rect 12887 7590 12899 7642
rect 12951 7590 12963 7642
rect 13015 7590 17146 7642
rect 17198 7590 17210 7642
rect 17262 7590 17274 7642
rect 17326 7590 17338 7642
rect 17390 7590 17402 7642
rect 17454 7590 18860 7642
rect 1104 7568 18860 7590
rect 382 7488 388 7540
rect 440 7528 446 7540
rect 440 7500 3556 7528
rect 440 7488 446 7500
rect 3418 7460 3424 7472
rect 3082 7432 3424 7460
rect 3418 7420 3424 7432
rect 3476 7420 3482 7472
rect 3528 7469 3556 7500
rect 3694 7488 3700 7540
rect 3752 7528 3758 7540
rect 9217 7531 9275 7537
rect 9217 7528 9229 7531
rect 3752 7500 9229 7528
rect 3752 7488 3758 7500
rect 9217 7497 9229 7500
rect 9263 7528 9275 7531
rect 9766 7528 9772 7540
rect 9263 7500 9772 7528
rect 9263 7497 9275 7500
rect 9217 7491 9275 7497
rect 9766 7488 9772 7500
rect 9824 7528 9830 7540
rect 9950 7528 9956 7540
rect 9824 7500 9956 7528
rect 9824 7488 9830 7500
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 10781 7531 10839 7537
rect 10152 7500 10732 7528
rect 3513 7463 3571 7469
rect 3513 7429 3525 7463
rect 3559 7460 3571 7463
rect 4065 7463 4123 7469
rect 4065 7460 4077 7463
rect 3559 7432 4077 7460
rect 3559 7429 3571 7432
rect 3513 7423 3571 7429
rect 4065 7429 4077 7432
rect 4111 7429 4123 7463
rect 4065 7423 4123 7429
rect 5810 7420 5816 7472
rect 5868 7460 5874 7472
rect 9582 7460 9588 7472
rect 5868 7432 9588 7460
rect 5868 7420 5874 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 1854 7352 1860 7404
rect 1912 7352 1918 7404
rect 5074 7352 5080 7404
rect 5132 7392 5138 7404
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 5132 7364 9965 7392
rect 5132 7352 5138 7364
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 1578 7284 1584 7336
rect 1636 7284 1642 7336
rect 1762 7284 1768 7336
rect 1820 7324 1826 7336
rect 2041 7327 2099 7333
rect 2041 7324 2053 7327
rect 1820 7296 2053 7324
rect 1820 7284 1826 7296
rect 2041 7293 2053 7296
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 3800 7327 3858 7333
rect 3800 7293 3812 7327
rect 3846 7324 3858 7327
rect 3846 7296 3924 7324
rect 3846 7293 3858 7296
rect 3800 7287 3858 7293
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3896 7188 3924 7296
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 10152 7324 10180 7500
rect 10502 7460 10508 7472
rect 10336 7432 10508 7460
rect 10336 7401 10364 7432
rect 10502 7420 10508 7432
rect 10560 7420 10566 7472
rect 10704 7460 10732 7500
rect 10781 7497 10793 7531
rect 10827 7528 10839 7531
rect 12618 7528 12624 7540
rect 10827 7500 12624 7528
rect 10827 7497 10839 7500
rect 10781 7491 10839 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 14182 7528 14188 7540
rect 13469 7500 14188 7528
rect 13469 7460 13497 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14366 7488 14372 7540
rect 14424 7488 14430 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15470 7528 15476 7540
rect 14783 7500 15476 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 16022 7528 16028 7540
rect 15896 7500 16028 7528
rect 15896 7488 15902 7500
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 17034 7488 17040 7540
rect 17092 7528 17098 7540
rect 17129 7531 17187 7537
rect 17129 7528 17141 7531
rect 17092 7500 17141 7528
rect 17092 7488 17098 7500
rect 17129 7497 17141 7500
rect 17175 7497 17187 7531
rect 17129 7491 17187 7497
rect 17494 7488 17500 7540
rect 17552 7488 17558 7540
rect 18230 7488 18236 7540
rect 18288 7528 18294 7540
rect 19242 7528 19248 7540
rect 18288 7500 19248 7528
rect 18288 7488 18294 7500
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 10704 7432 13497 7460
rect 15381 7463 15439 7469
rect 15381 7429 15393 7463
rect 15427 7460 15439 7463
rect 15746 7460 15752 7472
rect 15427 7432 15752 7460
rect 15427 7429 15439 7432
rect 10597 7419 10655 7425
rect 15381 7423 15439 7429
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 16298 7460 16304 7472
rect 15856 7432 16304 7460
rect 10597 7404 10609 7419
rect 10643 7404 10655 7419
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10594 7352 10600 7404
rect 10652 7352 10658 7404
rect 11146 7352 11152 7404
rect 11204 7352 11210 7404
rect 12158 7352 12164 7404
rect 12216 7352 12222 7404
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13504 7364 14289 7392
rect 13504 7352 13510 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 15010 7352 15016 7404
rect 15068 7392 15074 7404
rect 15856 7392 15884 7432
rect 16298 7420 16304 7432
rect 16356 7420 16362 7472
rect 16485 7463 16543 7469
rect 16485 7429 16497 7463
rect 16531 7460 16543 7463
rect 17954 7460 17960 7472
rect 16531 7432 17960 7460
rect 16531 7429 16543 7432
rect 16485 7423 16543 7429
rect 17954 7420 17960 7432
rect 18012 7420 18018 7472
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 15068 7364 15884 7392
rect 16040 7364 17049 7392
rect 15068 7352 15074 7364
rect 16040 7336 16068 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 17184 7364 18153 7392
rect 17184 7352 17190 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18325 7395 18383 7401
rect 18325 7361 18337 7395
rect 18371 7392 18383 7395
rect 18414 7392 18420 7404
rect 18371 7364 18420 7392
rect 18371 7361 18383 7364
rect 18325 7355 18383 7361
rect 18414 7352 18420 7364
rect 18472 7352 18478 7404
rect 9640 7296 10180 7324
rect 10505 7327 10563 7333
rect 9640 7284 9646 7296
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 13170 7324 13176 7336
rect 10551 7296 13176 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 14090 7284 14096 7336
rect 14148 7284 14154 7336
rect 16022 7284 16028 7336
rect 16080 7284 16086 7336
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7324 17003 7327
rect 17310 7324 17316 7336
rect 16991 7296 17316 7324
rect 16991 7293 17003 7296
rect 16945 7287 17003 7293
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 17402 7284 17408 7336
rect 17460 7324 17466 7336
rect 17681 7327 17739 7333
rect 17681 7324 17693 7327
rect 17460 7296 17693 7324
rect 17460 7284 17466 7296
rect 17681 7293 17693 7296
rect 17727 7293 17739 7327
rect 17681 7287 17739 7293
rect 17865 7327 17923 7333
rect 17865 7293 17877 7327
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 4798 7216 4804 7268
rect 4856 7256 4862 7268
rect 5445 7259 5503 7265
rect 5445 7256 5457 7259
rect 4856 7228 5457 7256
rect 4856 7216 4862 7228
rect 5445 7225 5457 7228
rect 5491 7256 5503 7259
rect 8294 7256 8300 7268
rect 5491 7228 8300 7256
rect 5491 7225 5503 7228
rect 5445 7219 5503 7225
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 10045 7259 10103 7265
rect 10045 7256 10057 7259
rect 10008 7228 10057 7256
rect 10008 7216 10014 7228
rect 10045 7225 10057 7228
rect 10091 7225 10103 7259
rect 10045 7219 10103 7225
rect 10520 7228 11468 7256
rect 3568 7160 3924 7188
rect 3568 7148 3574 7160
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10520 7188 10548 7228
rect 9824 7160 10548 7188
rect 11440 7188 11468 7228
rect 11514 7216 11520 7268
rect 11572 7256 11578 7268
rect 11974 7256 11980 7268
rect 11572 7228 11980 7256
rect 11572 7216 11578 7228
rect 11974 7216 11980 7228
rect 12032 7216 12038 7268
rect 12066 7216 12072 7268
rect 12124 7256 12130 7268
rect 12894 7256 12900 7268
rect 12124 7228 12900 7256
rect 12124 7216 12130 7228
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 13538 7216 13544 7268
rect 13596 7216 13602 7268
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 17880 7256 17908 7287
rect 17954 7284 17960 7336
rect 18012 7284 18018 7336
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7324 18107 7327
rect 18782 7324 18788 7336
rect 18095 7296 18788 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 13780 7228 17908 7256
rect 13780 7216 13786 7228
rect 13556 7188 13584 7216
rect 11440 7160 13584 7188
rect 9824 7148 9830 7160
rect 13630 7148 13636 7200
rect 13688 7148 13694 7200
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 18064 7188 18092 7287
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 15795 7160 18092 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 2133 6987 2191 6993
rect 2133 6953 2145 6987
rect 2179 6984 2191 6987
rect 2314 6984 2320 6996
rect 2179 6956 2320 6984
rect 2179 6953 2191 6956
rect 2133 6947 2191 6953
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7113 6987 7171 6993
rect 7113 6984 7125 6987
rect 6972 6956 7125 6984
rect 6972 6944 6978 6956
rect 7113 6953 7125 6956
rect 7159 6953 7171 6987
rect 7113 6947 7171 6953
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6984 9919 6987
rect 10502 6984 10508 6996
rect 9907 6956 10508 6984
rect 9907 6953 9919 6956
rect 9861 6947 9919 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 11897 6987 11955 6993
rect 11897 6984 11909 6987
rect 11756 6956 11909 6984
rect 11756 6944 11762 6956
rect 11897 6953 11909 6956
rect 11943 6953 11955 6987
rect 11897 6947 11955 6953
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 12986 6984 12992 6996
rect 12216 6956 12992 6984
rect 12216 6944 12222 6956
rect 12986 6944 12992 6956
rect 13044 6984 13050 6996
rect 13354 6984 13360 6996
rect 13044 6956 13360 6984
rect 13044 6944 13050 6956
rect 13354 6944 13360 6956
rect 13412 6984 13418 6996
rect 14277 6987 14335 6993
rect 14277 6984 14289 6987
rect 13412 6956 14289 6984
rect 13412 6944 13418 6956
rect 14277 6953 14289 6956
rect 14323 6953 14335 6987
rect 14277 6947 14335 6953
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 16298 6984 16304 6996
rect 15620 6956 16304 6984
rect 15620 6944 15626 6956
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 16669 6987 16727 6993
rect 16669 6953 16681 6987
rect 16715 6984 16727 6987
rect 17310 6984 17316 6996
rect 16715 6956 17316 6984
rect 16715 6953 16727 6956
rect 16669 6947 16727 6953
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 1762 6876 1768 6928
rect 1820 6916 1826 6928
rect 2593 6919 2651 6925
rect 2593 6916 2605 6919
rect 1820 6888 2605 6916
rect 1820 6876 1826 6888
rect 2593 6885 2605 6888
rect 2639 6916 2651 6919
rect 2682 6916 2688 6928
rect 2639 6888 2688 6916
rect 2639 6885 2651 6888
rect 2593 6879 2651 6885
rect 2682 6876 2688 6888
rect 2740 6916 2746 6928
rect 2740 6888 3648 6916
rect 2740 6876 2746 6888
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 3620 6848 3648 6888
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 10413 6919 10471 6925
rect 10413 6916 10425 6919
rect 8352 6888 10425 6916
rect 8352 6876 8358 6888
rect 10413 6885 10425 6888
rect 10459 6885 10471 6919
rect 10413 6879 10471 6885
rect 12710 6876 12716 6928
rect 12768 6876 12774 6928
rect 12894 6876 12900 6928
rect 12952 6916 12958 6928
rect 13722 6916 13728 6928
rect 12952 6888 13728 6916
rect 12952 6876 12958 6888
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 15930 6876 15936 6928
rect 15988 6916 15994 6928
rect 17865 6919 17923 6925
rect 17865 6916 17877 6919
rect 15988 6888 17877 6916
rect 15988 6876 15994 6888
rect 17865 6885 17877 6888
rect 17911 6885 17923 6919
rect 17865 6879 17923 6885
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 1452 6820 3096 6848
rect 3620 6820 4445 6848
rect 1452 6808 1458 6820
rect 1854 6740 1860 6792
rect 1912 6740 1918 6792
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2314 6780 2320 6792
rect 1995 6752 2320 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 2774 6740 2780 6792
rect 2832 6740 2838 6792
rect 2958 6740 2964 6792
rect 3016 6740 3022 6792
rect 3068 6780 3096 6820
rect 4433 6817 4445 6820
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 8389 6851 8447 6857
rect 8389 6848 8401 6851
rect 6788 6820 8401 6848
rect 6788 6808 6794 6820
rect 8389 6817 8401 6820
rect 8435 6817 8447 6851
rect 8389 6811 8447 6817
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 9364 6820 12173 6848
rect 9364 6808 9370 6820
rect 12161 6817 12173 6820
rect 12207 6848 12219 6851
rect 13630 6848 13636 6860
rect 12207 6820 13636 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 17586 6848 17592 6860
rect 16448 6820 17592 6848
rect 16448 6808 16454 6820
rect 17586 6808 17592 6820
rect 17644 6848 17650 6860
rect 17644 6820 17816 6848
rect 17644 6808 17650 6820
rect 3068 6752 4200 6780
rect 2130 6672 2136 6724
rect 2188 6712 2194 6724
rect 2498 6712 2504 6724
rect 2188 6684 2504 6712
rect 2188 6672 2194 6684
rect 2498 6672 2504 6684
rect 2556 6672 2562 6724
rect 2976 6712 3004 6740
rect 2792 6684 3004 6712
rect 3513 6715 3571 6721
rect 2792 6656 2820 6684
rect 3513 6681 3525 6715
rect 3559 6681 3571 6715
rect 3513 6675 3571 6681
rect 1670 6604 1676 6656
rect 1728 6604 1734 6656
rect 2774 6604 2780 6656
rect 2832 6604 2838 6656
rect 2958 6604 2964 6656
rect 3016 6604 3022 6656
rect 3418 6604 3424 6656
rect 3476 6604 3482 6656
rect 3528 6644 3556 6675
rect 3602 6672 3608 6724
rect 3660 6712 3666 6724
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3660 6684 3801 6712
rect 3660 6672 3666 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 4062 6672 4068 6724
rect 4120 6672 4126 6724
rect 4172 6712 4200 6752
rect 4338 6740 4344 6792
rect 4396 6740 4402 6792
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 8573 6783 8631 6789
rect 8573 6780 8585 6783
rect 8343 6752 8585 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 8573 6749 8585 6752
rect 8619 6780 8631 6783
rect 8662 6780 8668 6792
rect 8619 6752 8668 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 5353 6715 5411 6721
rect 5353 6712 5365 6715
rect 4172 6684 5365 6712
rect 5353 6681 5365 6684
rect 5399 6681 5411 6715
rect 5353 6675 5411 6681
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 5684 6684 5934 6712
rect 5684 6672 5690 6684
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7392 6712 7420 6743
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 10778 6740 10784 6792
rect 10836 6740 10842 6792
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12584 6752 12909 6780
rect 12584 6740 12590 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 7248 6684 7420 6712
rect 7484 6684 10640 6712
rect 7248 6672 7254 6684
rect 3694 6644 3700 6656
rect 3528 6616 3700 6644
rect 3694 6604 3700 6616
rect 3752 6644 3758 6656
rect 7484 6644 7512 6684
rect 3752 6616 7512 6644
rect 8757 6647 8815 6653
rect 3752 6604 3758 6616
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 9582 6644 9588 6656
rect 8803 6616 9588 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 10612 6644 10640 6684
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 12158 6712 12164 6724
rect 11848 6684 12164 6712
rect 11848 6672 11854 6684
rect 12158 6672 12164 6684
rect 12216 6672 12222 6724
rect 12250 6672 12256 6724
rect 12308 6672 12314 6724
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 12621 6715 12679 6721
rect 12621 6712 12633 6715
rect 12400 6684 12633 6712
rect 12400 6672 12406 6684
rect 12621 6681 12633 6684
rect 12667 6712 12679 6715
rect 12912 6712 12940 6743
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13081 6783 13139 6789
rect 13081 6780 13093 6783
rect 13044 6752 13093 6780
rect 13044 6740 13050 6752
rect 13081 6749 13093 6752
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 14148 6752 17417 6780
rect 14148 6740 14154 6752
rect 17405 6749 17417 6752
rect 17451 6780 17463 6783
rect 17678 6780 17684 6792
rect 17451 6752 17684 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 17788 6789 17816 6820
rect 17773 6783 17831 6789
rect 17773 6749 17785 6783
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 18104 6752 18337 6780
rect 18104 6740 18110 6752
rect 18325 6749 18337 6752
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 13725 6715 13783 6721
rect 13725 6712 13737 6715
rect 12667 6684 12848 6712
rect 12912 6684 13737 6712
rect 12667 6681 12679 6684
rect 12621 6675 12679 6681
rect 11054 6644 11060 6656
rect 10612 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 12710 6644 12716 6656
rect 11296 6616 12716 6644
rect 11296 6604 11302 6616
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 12820 6644 12848 6684
rect 13725 6681 13737 6684
rect 13771 6681 13783 6715
rect 13725 6675 13783 6681
rect 16850 6672 16856 6724
rect 16908 6712 16914 6724
rect 17310 6712 17316 6724
rect 16908 6684 17316 6712
rect 16908 6672 16914 6684
rect 17310 6672 17316 6684
rect 17368 6672 17374 6724
rect 13814 6644 13820 6656
rect 12820 6616 13820 6644
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 16942 6604 16948 6656
rect 17000 6604 17006 6656
rect 1104 6554 18860 6576
rect 1104 6502 3829 6554
rect 3881 6502 3893 6554
rect 3945 6502 3957 6554
rect 4009 6502 4021 6554
rect 4073 6502 4085 6554
rect 4137 6502 8268 6554
rect 8320 6502 8332 6554
rect 8384 6502 8396 6554
rect 8448 6502 8460 6554
rect 8512 6502 8524 6554
rect 8576 6502 12707 6554
rect 12759 6502 12771 6554
rect 12823 6502 12835 6554
rect 12887 6502 12899 6554
rect 12951 6502 12963 6554
rect 13015 6502 17146 6554
rect 17198 6502 17210 6554
rect 17262 6502 17274 6554
rect 17326 6502 17338 6554
rect 17390 6502 17402 6554
rect 17454 6502 18860 6554
rect 1104 6480 18860 6502
rect 3237 6443 3295 6449
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 5166 6440 5172 6452
rect 3283 6412 5172 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 6546 6440 6552 6452
rect 5307 6412 6552 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 1118 6332 1124 6384
rect 1176 6372 1182 6384
rect 1176 6344 1992 6372
rect 1176 6332 1182 6344
rect 1394 6264 1400 6316
rect 1452 6304 1458 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1452 6276 1869 6304
rect 1452 6264 1458 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 1964 6304 1992 6344
rect 2314 6332 2320 6384
rect 2372 6372 2378 6384
rect 2409 6375 2467 6381
rect 2409 6372 2421 6375
rect 2372 6344 2421 6372
rect 2372 6332 2378 6344
rect 2409 6341 2421 6344
rect 2455 6372 2467 6375
rect 4522 6372 4528 6384
rect 2455 6344 4528 6372
rect 2455 6341 2467 6344
rect 2409 6335 2467 6341
rect 4522 6332 4528 6344
rect 4580 6332 4586 6384
rect 5537 6375 5595 6381
rect 5537 6372 5549 6375
rect 5092 6344 5549 6372
rect 2869 6307 2927 6313
rect 2869 6304 2881 6307
rect 1964 6276 2881 6304
rect 1857 6267 1915 6273
rect 2869 6273 2881 6276
rect 2915 6304 2927 6307
rect 4154 6304 4160 6316
rect 2915 6276 4160 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 842 6196 848 6248
rect 900 6236 906 6248
rect 1581 6239 1639 6245
rect 1581 6236 1593 6239
rect 900 6208 1593 6236
rect 900 6196 906 6208
rect 1581 6205 1593 6208
rect 1627 6205 1639 6239
rect 1581 6199 1639 6205
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6205 2743 6239
rect 2685 6199 2743 6205
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 2823 6208 4108 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 2700 6168 2728 6199
rect 2866 6168 2872 6180
rect 2700 6140 2872 6168
rect 2866 6128 2872 6140
rect 2924 6128 2930 6180
rect 3694 6128 3700 6180
rect 3752 6128 3758 6180
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 2958 6100 2964 6112
rect 1912 6072 2964 6100
rect 1912 6060 1918 6072
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 4080 6100 4108 6208
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4801 6239 4859 6245
rect 4801 6236 4813 6239
rect 4304 6208 4813 6236
rect 4304 6196 4310 6208
rect 4801 6205 4813 6208
rect 4847 6236 4859 6239
rect 5092 6236 5120 6344
rect 5537 6341 5549 6344
rect 5583 6341 5595 6375
rect 5537 6335 5595 6341
rect 5626 6332 5632 6384
rect 5684 6332 5690 6384
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5741 6313 5769 6412
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 6638 6400 6644 6452
rect 6696 6400 6702 6452
rect 6730 6400 6736 6452
rect 6788 6400 6794 6452
rect 7098 6400 7104 6452
rect 7156 6400 7162 6452
rect 8386 6440 8392 6452
rect 7208 6412 8392 6440
rect 7208 6372 7236 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 9456 6412 9689 6440
rect 9456 6400 9462 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 9677 6403 9735 6409
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 11238 6440 11244 6452
rect 10192 6412 11244 6440
rect 10192 6400 10198 6412
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 11480 6412 12265 6440
rect 11480 6400 11486 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 13078 6440 13084 6452
rect 12253 6403 12311 6409
rect 12544 6412 13084 6440
rect 6104 6344 7236 6372
rect 5373 6307 5431 6313
rect 5373 6304 5385 6307
rect 5224 6276 5385 6304
rect 5224 6264 5230 6276
rect 5368 6273 5385 6276
rect 5419 6273 5431 6307
rect 5368 6267 5431 6273
rect 5726 6307 5784 6313
rect 5726 6273 5738 6307
rect 5772 6273 5784 6307
rect 5726 6267 5784 6273
rect 4847 6208 5120 6236
rect 5368 6236 5396 6267
rect 5810 6236 5816 6248
rect 5368 6208 5816 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 4157 6171 4215 6177
rect 4157 6137 4169 6171
rect 4203 6168 4215 6171
rect 4338 6168 4344 6180
rect 4203 6140 4344 6168
rect 4203 6137 4215 6140
rect 4157 6131 4215 6137
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 4890 6128 4896 6180
rect 4948 6128 4954 6180
rect 5905 6171 5963 6177
rect 5905 6137 5917 6171
rect 5951 6168 5963 6171
rect 5994 6168 6000 6180
rect 5951 6140 6000 6168
rect 5951 6137 5963 6140
rect 5905 6131 5963 6137
rect 5994 6128 6000 6140
rect 6052 6128 6058 6180
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 4080 6072 4537 6100
rect 4525 6069 4537 6072
rect 4571 6100 4583 6103
rect 4908 6100 4936 6128
rect 6104 6100 6132 6344
rect 8110 6332 8116 6384
rect 8168 6332 8174 6384
rect 9122 6332 9128 6384
rect 9180 6332 9186 6384
rect 9324 6372 9352 6400
rect 9324 6344 9444 6372
rect 9416 6313 9444 6344
rect 9490 6332 9496 6384
rect 9548 6332 9554 6384
rect 10042 6332 10048 6384
rect 10100 6332 10106 6384
rect 12544 6372 12572 6412
rect 13078 6400 13084 6412
rect 13136 6440 13142 6452
rect 13541 6443 13599 6449
rect 13541 6440 13553 6443
rect 13136 6412 13553 6440
rect 13136 6400 13142 6412
rect 13541 6409 13553 6412
rect 13587 6440 13599 6443
rect 14734 6440 14740 6452
rect 13587 6412 14740 6440
rect 13587 6409 13599 6412
rect 13541 6403 13599 6409
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 17034 6400 17040 6452
rect 17092 6400 17098 6452
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17770 6440 17776 6452
rect 17543 6412 17776 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 17865 6443 17923 6449
rect 17865 6409 17877 6443
rect 17911 6440 17923 6443
rect 18506 6440 18512 6452
rect 17911 6412 18512 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 11808 6344 12572 6372
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9766 6304 9772 6316
rect 9447 6276 9772 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10594 6304 10600 6316
rect 10459 6276 10600 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10594 6264 10600 6276
rect 10652 6304 10658 6316
rect 11514 6304 11520 6316
rect 10652 6276 11520 6304
rect 10652 6264 10658 6276
rect 11514 6264 11520 6276
rect 11572 6264 11578 6316
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 7466 6236 7472 6248
rect 6604 6208 7472 6236
rect 6604 6196 6610 6208
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 11808 6236 11836 6344
rect 12618 6332 12624 6384
rect 12676 6372 12682 6384
rect 12897 6375 12955 6381
rect 12897 6372 12909 6375
rect 12676 6344 12909 6372
rect 12676 6332 12682 6344
rect 12897 6341 12909 6344
rect 12943 6341 12955 6375
rect 12897 6335 12955 6341
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 11940 6276 12449 6304
rect 11940 6264 11946 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 12526 6264 12532 6316
rect 12584 6264 12590 6316
rect 13078 6264 13084 6316
rect 13136 6264 13142 6316
rect 13265 6307 13323 6313
rect 13265 6304 13277 6307
rect 13188 6276 13277 6304
rect 8812 6208 11836 6236
rect 8812 6196 8818 6208
rect 12802 6196 12808 6248
rect 12860 6196 12866 6248
rect 12986 6196 12992 6248
rect 13044 6236 13050 6248
rect 13188 6236 13216 6276
rect 13265 6273 13277 6276
rect 13311 6304 13323 6307
rect 13998 6304 14004 6316
rect 13311 6276 14004 6304
rect 13311 6273 13323 6276
rect 13265 6267 13323 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 13044 6208 13216 6236
rect 13044 6196 13050 6208
rect 6914 6128 6920 6180
rect 6972 6168 6978 6180
rect 6972 6140 7512 6168
rect 6972 6128 6978 6140
rect 4571 6072 6132 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 7377 6103 7435 6109
rect 7377 6100 7389 6103
rect 6880 6072 7389 6100
rect 6880 6060 6886 6072
rect 7377 6069 7389 6072
rect 7423 6069 7435 6103
rect 7484 6100 7512 6140
rect 7650 6128 7656 6180
rect 7708 6168 7714 6180
rect 8110 6168 8116 6180
rect 7708 6140 8116 6168
rect 7708 6128 7714 6140
rect 8110 6128 8116 6140
rect 8168 6128 8174 6180
rect 10134 6168 10140 6180
rect 9324 6140 10140 6168
rect 9324 6100 9352 6140
rect 10134 6128 10140 6140
rect 10192 6168 10198 6180
rect 11977 6171 12035 6177
rect 11977 6168 11989 6171
rect 10192 6140 11989 6168
rect 10192 6128 10198 6140
rect 11977 6137 11989 6140
rect 12023 6137 12035 6171
rect 11977 6131 12035 6137
rect 7484 6072 9352 6100
rect 11992 6100 12020 6131
rect 12066 6128 12072 6180
rect 12124 6168 12130 6180
rect 16022 6168 16028 6180
rect 12124 6140 16028 6168
rect 12124 6128 12130 6140
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 12713 6103 12771 6109
rect 12713 6100 12725 6103
rect 11992 6072 12725 6100
rect 7377 6063 7435 6069
rect 12713 6069 12725 6072
rect 12759 6100 12771 6103
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 12759 6072 18245 6100
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 18233 6069 18245 6072
rect 18279 6100 18291 6103
rect 18414 6100 18420 6112
rect 18279 6072 18420 6100
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 2133 5899 2191 5905
rect 2133 5865 2145 5899
rect 2179 5896 2191 5899
rect 2222 5896 2228 5908
rect 2179 5868 2228 5896
rect 2179 5865 2191 5868
rect 2133 5859 2191 5865
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 2593 5899 2651 5905
rect 2593 5896 2605 5899
rect 2556 5868 2605 5896
rect 2556 5856 2562 5868
rect 2593 5865 2605 5868
rect 2639 5865 2651 5899
rect 2593 5859 2651 5865
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 2924 5868 3985 5896
rect 2924 5856 2930 5868
rect 3973 5865 3985 5868
rect 4019 5865 4031 5899
rect 3973 5859 4031 5865
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 4764 5868 5365 5896
rect 4764 5856 4770 5868
rect 5353 5865 5365 5868
rect 5399 5896 5411 5899
rect 5994 5896 6000 5908
rect 5399 5868 6000 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 6270 5856 6276 5908
rect 6328 5856 6334 5908
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 7745 5899 7803 5905
rect 7745 5896 7757 5899
rect 6512 5868 7757 5896
rect 6512 5856 6518 5868
rect 7745 5865 7757 5868
rect 7791 5865 7803 5899
rect 7745 5859 7803 5865
rect 2038 5828 2044 5840
rect 1872 5800 2044 5828
rect 1872 5701 1900 5800
rect 2038 5788 2044 5800
rect 2096 5788 2102 5840
rect 7101 5831 7159 5837
rect 7101 5797 7113 5831
rect 7147 5797 7159 5831
rect 7101 5791 7159 5797
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2406 5760 2412 5772
rect 2271 5732 2412 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 2958 5720 2964 5772
rect 3016 5760 3022 5772
rect 3016 5732 6224 5760
rect 3016 5720 3022 5732
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1946 5652 1952 5704
rect 2004 5652 2010 5704
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2314 5692 2320 5704
rect 2087 5664 2320 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5592 5664 5917 5692
rect 5592 5652 5598 5664
rect 5905 5661 5917 5664
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 6052 5664 6101 5692
rect 6052 5652 6058 5664
rect 6089 5661 6101 5664
rect 6135 5661 6147 5695
rect 6196 5692 6224 5732
rect 6362 5720 6368 5772
rect 6420 5760 6426 5772
rect 6457 5763 6515 5769
rect 6457 5760 6469 5763
rect 6420 5732 6469 5760
rect 6420 5720 6426 5732
rect 6457 5729 6469 5732
rect 6503 5729 6515 5763
rect 6457 5723 6515 5729
rect 7116 5692 7144 5791
rect 7760 5760 7788 5859
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 12526 5896 12532 5908
rect 8444 5868 12532 5896
rect 8444 5856 8450 5868
rect 12526 5856 12532 5868
rect 12584 5896 12590 5908
rect 13538 5896 13544 5908
rect 12584 5868 13544 5896
rect 12584 5856 12590 5868
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14182 5856 14188 5908
rect 14240 5856 14246 5908
rect 16850 5896 16856 5908
rect 14292 5868 16856 5896
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 10318 5828 10324 5840
rect 8536 5800 10324 5828
rect 8536 5788 8542 5800
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 11204 5800 12572 5828
rect 11204 5788 11210 5800
rect 7760 5758 8156 5760
rect 7760 5732 8248 5758
rect 8128 5730 8248 5732
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 6196 5664 6776 5692
rect 7116 5664 8125 5692
rect 6089 5655 6147 5661
rect 1578 5584 1584 5636
rect 1636 5584 1642 5636
rect 3605 5627 3663 5633
rect 3605 5593 3617 5627
rect 3651 5624 3663 5627
rect 4154 5624 4160 5636
rect 3651 5596 4160 5624
rect 3651 5593 3663 5596
rect 3605 5587 3663 5593
rect 4154 5584 4160 5596
rect 4212 5624 4218 5636
rect 5166 5624 5172 5636
rect 4212 5596 5172 5624
rect 4212 5584 4218 5596
rect 5166 5584 5172 5596
rect 5224 5584 5230 5636
rect 6454 5584 6460 5636
rect 6512 5624 6518 5636
rect 6641 5627 6699 5633
rect 6641 5624 6653 5627
rect 6512 5596 6653 5624
rect 6512 5584 6518 5596
rect 6641 5593 6653 5596
rect 6687 5593 6699 5627
rect 6748 5624 6776 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8220 5692 8248 5730
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 10226 5760 10232 5772
rect 8628 5732 10232 5760
rect 8628 5720 8634 5732
rect 10226 5720 10232 5732
rect 10284 5760 10290 5772
rect 10686 5760 10692 5772
rect 10284 5732 10692 5760
rect 10284 5720 10290 5732
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 9950 5692 9956 5704
rect 8220 5664 9956 5692
rect 8113 5655 8171 5661
rect 9950 5652 9956 5664
rect 10008 5692 10014 5704
rect 11882 5692 11888 5704
rect 10008 5664 11888 5692
rect 10008 5652 10014 5664
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 12544 5692 12572 5800
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 14292 5828 14320 5868
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17586 5856 17592 5908
rect 17644 5856 17650 5908
rect 18049 5899 18107 5905
rect 18049 5865 18061 5899
rect 18095 5896 18107 5899
rect 18414 5896 18420 5908
rect 18095 5868 18420 5896
rect 18095 5865 18107 5868
rect 18049 5859 18107 5865
rect 18414 5856 18420 5868
rect 18472 5896 18478 5908
rect 18874 5896 18880 5908
rect 18472 5868 18880 5896
rect 18472 5856 18478 5868
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 12676 5800 14320 5828
rect 12676 5788 12682 5800
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 12860 5732 12909 5760
rect 12860 5720 12866 5732
rect 12897 5729 12909 5732
rect 12943 5760 12955 5763
rect 13078 5760 13084 5772
rect 12943 5732 13084 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 13630 5720 13636 5772
rect 13688 5760 13694 5772
rect 15933 5763 15991 5769
rect 15933 5760 15945 5763
rect 13688 5732 15945 5760
rect 13688 5720 13694 5732
rect 15933 5729 15945 5732
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 18104 5732 18429 5760
rect 18104 5720 18110 5732
rect 18417 5729 18429 5732
rect 18463 5729 18475 5763
rect 18417 5723 18475 5729
rect 13998 5692 14004 5704
rect 12544 5664 14004 5692
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 8018 5624 8024 5636
rect 6748 5596 8024 5624
rect 6641 5587 6699 5593
rect 8018 5584 8024 5596
rect 8076 5584 8082 5636
rect 8309 5627 8367 5633
rect 8309 5593 8321 5627
rect 8355 5624 8367 5627
rect 8478 5624 8484 5636
rect 8355 5596 8484 5624
rect 8355 5593 8367 5596
rect 8309 5587 8367 5593
rect 8478 5584 8484 5596
rect 8536 5584 8542 5636
rect 9398 5584 9404 5636
rect 9456 5584 9462 5636
rect 10594 5624 10600 5636
rect 9646 5596 10600 5624
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 5074 5556 5080 5568
rect 2924 5528 5080 5556
rect 2924 5516 2930 5528
rect 5074 5516 5080 5528
rect 5132 5556 5138 5568
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 5132 5528 5733 5556
rect 5132 5516 5138 5528
rect 5721 5525 5733 5528
rect 5767 5525 5779 5559
rect 5721 5519 5779 5525
rect 5902 5516 5908 5568
rect 5960 5556 5966 5568
rect 6730 5556 6736 5568
rect 5960 5528 6736 5556
rect 5960 5516 5966 5528
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 9646 5556 9674 5596
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 11238 5584 11244 5636
rect 11296 5624 11302 5636
rect 14090 5624 14096 5636
rect 11296 5596 14096 5624
rect 11296 5584 11302 5596
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 15102 5584 15108 5636
rect 15160 5584 15166 5636
rect 15657 5627 15715 5633
rect 15657 5593 15669 5627
rect 15703 5593 15715 5627
rect 15657 5587 15715 5593
rect 7524 5528 9674 5556
rect 7524 5516 7530 5528
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 11756 5528 12541 5556
rect 11756 5516 11762 5528
rect 12529 5525 12541 5528
rect 12575 5556 12587 5559
rect 12986 5556 12992 5568
rect 12575 5528 12992 5556
rect 12575 5525 12587 5528
rect 12529 5519 12587 5525
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 15672 5556 15700 5587
rect 13964 5528 15700 5556
rect 13964 5516 13970 5528
rect 1104 5466 18860 5488
rect 1104 5414 3829 5466
rect 3881 5414 3893 5466
rect 3945 5414 3957 5466
rect 4009 5414 4021 5466
rect 4073 5414 4085 5466
rect 4137 5414 8268 5466
rect 8320 5414 8332 5466
rect 8384 5414 8396 5466
rect 8448 5414 8460 5466
rect 8512 5414 8524 5466
rect 8576 5414 12707 5466
rect 12759 5414 12771 5466
rect 12823 5414 12835 5466
rect 12887 5414 12899 5466
rect 12951 5414 12963 5466
rect 13015 5414 17146 5466
rect 17198 5414 17210 5466
rect 17262 5414 17274 5466
rect 17326 5414 17338 5466
rect 17390 5414 17402 5466
rect 17454 5414 18860 5466
rect 1104 5392 18860 5414
rect 2314 5312 2320 5364
rect 2372 5312 2378 5364
rect 4154 5352 4160 5364
rect 3068 5324 4160 5352
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 2590 5216 2596 5228
rect 1903 5188 2596 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2866 5216 2872 5228
rect 2731 5188 2872 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 2958 5176 2964 5228
rect 3016 5176 3022 5228
rect 842 5108 848 5160
rect 900 5148 906 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 900 5120 1593 5148
rect 900 5108 906 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 3068 5148 3096 5324
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 9214 5352 9220 5364
rect 4304 5324 9220 5352
rect 4304 5312 4310 5324
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9456 5324 10057 5352
rect 9456 5312 9462 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10045 5315 10103 5321
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18141 5355 18199 5361
rect 18141 5352 18153 5355
rect 18012 5324 18153 5352
rect 18012 5312 18018 5324
rect 18141 5321 18153 5324
rect 18187 5321 18199 5355
rect 18141 5315 18199 5321
rect 4798 5284 4804 5296
rect 4738 5256 4804 5284
rect 4798 5244 4804 5256
rect 4856 5284 4862 5296
rect 7006 5284 7012 5296
rect 4856 5256 7012 5284
rect 4856 5244 4862 5256
rect 7006 5244 7012 5256
rect 7064 5284 7070 5296
rect 9493 5287 9551 5293
rect 7064 5256 8326 5284
rect 7064 5244 7070 5256
rect 9493 5253 9505 5287
rect 9539 5284 9551 5287
rect 15654 5284 15660 5296
rect 9539 5256 15660 5284
rect 9539 5253 9551 5256
rect 9493 5247 9551 5253
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 18690 5284 18696 5296
rect 15764 5256 18696 5284
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 5776 5188 6561 5216
rect 5776 5176 5782 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 6788 5188 7389 5216
rect 6788 5176 6794 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 2823 5120 3096 5148
rect 3237 5151 3295 5157
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 3513 5151 3571 5157
rect 3283 5120 3372 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3344 5012 3372 5120
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 3559 5120 5457 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 5445 5117 5457 5120
rect 5491 5148 5503 5151
rect 6638 5148 6644 5160
rect 5491 5120 6644 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 7392 5148 7420 5179
rect 9766 5176 9772 5228
rect 9824 5176 9830 5228
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 7392 5120 7972 5148
rect 5350 5080 5356 5092
rect 4540 5052 5356 5080
rect 3510 5012 3516 5024
rect 3344 4984 3516 5012
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4540 5012 4568 5052
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 4212 4984 4568 5012
rect 4212 4972 4218 4984
rect 4982 4972 4988 5024
rect 5040 4972 5046 5024
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 6546 5012 6552 5024
rect 6420 4984 6552 5012
rect 6420 4972 6426 4984
rect 6546 4972 6552 4984
rect 6604 5012 6610 5024
rect 7745 5015 7803 5021
rect 7745 5012 7757 5015
rect 6604 4984 7757 5012
rect 6604 4972 6610 4984
rect 7745 4981 7757 4984
rect 7791 4981 7803 5015
rect 7944 5012 7972 5120
rect 8018 5108 8024 5160
rect 8076 5108 8082 5160
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 15764 5148 15792 5256
rect 18690 5244 18696 5256
rect 18748 5244 18754 5296
rect 18322 5176 18328 5228
rect 18380 5176 18386 5228
rect 18414 5176 18420 5228
rect 18472 5176 18478 5228
rect 8536 5120 15792 5148
rect 8536 5108 8542 5120
rect 16298 5108 16304 5160
rect 16356 5148 16362 5160
rect 17773 5151 17831 5157
rect 17773 5148 17785 5151
rect 16356 5120 17785 5148
rect 16356 5108 16362 5120
rect 17773 5117 17785 5120
rect 17819 5148 17831 5151
rect 18141 5151 18199 5157
rect 18141 5148 18153 5151
rect 17819 5120 18153 5148
rect 17819 5117 17831 5120
rect 17773 5111 17831 5117
rect 18141 5117 18153 5120
rect 18187 5117 18199 5151
rect 18141 5111 18199 5117
rect 17862 5080 17868 5092
rect 9692 5052 17868 5080
rect 9692 5012 9720 5052
rect 17862 5040 17868 5052
rect 17920 5040 17926 5092
rect 7944 4984 9720 5012
rect 7745 4975 7803 4981
rect 14826 4972 14832 5024
rect 14884 5012 14890 5024
rect 18046 5012 18052 5024
rect 14884 4984 18052 5012
rect 14884 4972 14890 4984
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 2038 4768 2044 4820
rect 2096 4808 2102 4820
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 2096 4780 2145 4808
rect 2096 4768 2102 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 2133 4771 2191 4777
rect 2590 4768 2596 4820
rect 2648 4768 2654 4820
rect 2958 4768 2964 4820
rect 3016 4808 3022 4820
rect 3145 4811 3203 4817
rect 3145 4808 3157 4811
rect 3016 4780 3157 4808
rect 3016 4768 3022 4780
rect 3145 4777 3157 4780
rect 3191 4808 3203 4811
rect 4154 4808 4160 4820
rect 3191 4780 4160 4808
rect 3191 4777 3203 4780
rect 3145 4771 3203 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5040 4780 13124 4808
rect 5040 4768 5046 4780
rect 2866 4700 2872 4752
rect 2924 4740 2930 4752
rect 3421 4743 3479 4749
rect 3421 4740 3433 4743
rect 2924 4712 3433 4740
rect 2924 4700 2930 4712
rect 3421 4709 3433 4712
rect 3467 4709 3479 4743
rect 3421 4703 3479 4709
rect 3878 4700 3884 4752
rect 3936 4740 3942 4752
rect 4617 4743 4675 4749
rect 4617 4740 4629 4743
rect 3936 4712 4629 4740
rect 3936 4700 3942 4712
rect 4617 4709 4629 4712
rect 4663 4709 4675 4743
rect 6089 4743 6147 4749
rect 6089 4740 6101 4743
rect 4617 4703 4675 4709
rect 5276 4712 6101 4740
rect 5276 4681 5304 4712
rect 6089 4709 6101 4712
rect 6135 4740 6147 4743
rect 6454 4740 6460 4752
rect 6135 4712 6460 4740
rect 6135 4709 6147 4712
rect 6089 4703 6147 4709
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 6638 4700 6644 4752
rect 6696 4740 6702 4752
rect 8478 4740 8484 4752
rect 6696 4712 8484 4740
rect 6696 4700 6702 4712
rect 8478 4700 8484 4712
rect 8536 4700 8542 4752
rect 13096 4740 13124 4780
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 13228 4780 14197 4808
rect 13228 4768 13234 4780
rect 14185 4777 14197 4780
rect 14231 4777 14243 4811
rect 14185 4771 14243 4777
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 14826 4808 14832 4820
rect 14691 4780 14832 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 14366 4740 14372 4752
rect 12406 4712 13032 4740
rect 13096 4712 14372 4740
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4672 4215 4675
rect 5261 4675 5319 4681
rect 4203 4644 5028 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 5000 4616 5028 4644
rect 5261 4641 5273 4675
rect 5307 4641 5319 4675
rect 5261 4635 5319 4641
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 8757 4675 8815 4681
rect 7340 4644 7498 4672
rect 7340 4632 7346 4644
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9674 4672 9680 4684
rect 8803 4644 9680 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 1854 4564 1860 4616
rect 1912 4564 1918 4616
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4798 4604 4804 4616
rect 4396 4576 4804 4604
rect 4396 4564 4402 4576
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 4982 4564 4988 4616
rect 5040 4564 5046 4616
rect 7558 4564 7564 4616
rect 7616 4564 7622 4616
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 12406 4604 12434 4712
rect 13004 4672 13032 4712
rect 14366 4700 14372 4712
rect 14424 4700 14430 4752
rect 13909 4675 13967 4681
rect 13004 4644 13676 4672
rect 8435 4576 12434 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 13648 4548 13676 4644
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 14090 4672 14096 4684
rect 13955 4644 14096 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 14660 4672 14688 4771
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 17037 4743 17095 4749
rect 17037 4709 17049 4743
rect 17083 4740 17095 4743
rect 19150 4740 19156 4752
rect 17083 4712 19156 4740
rect 17083 4709 17095 4712
rect 17037 4703 17095 4709
rect 19150 4700 19156 4712
rect 19208 4700 19214 4752
rect 14292 4644 14688 4672
rect 14292 4613 14320 4644
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 16908 4644 17264 4672
rect 16908 4632 16914 4644
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 17236 4613 17264 4644
rect 17221 4607 17279 4613
rect 14516 4576 16252 4604
rect 14516 4564 14522 4576
rect 842 4496 848 4548
rect 900 4536 906 4548
rect 1581 4539 1639 4545
rect 1581 4536 1593 4539
rect 900 4508 1593 4536
rect 900 4496 906 4508
rect 1581 4505 1593 4508
rect 1627 4505 1639 4539
rect 1581 4499 1639 4505
rect 3326 4496 3332 4548
rect 3384 4536 3390 4548
rect 13078 4536 13084 4548
rect 3384 4508 13084 4536
rect 3384 4496 3390 4508
rect 13078 4496 13084 4508
rect 13136 4496 13142 4548
rect 13630 4496 13636 4548
rect 13688 4536 13694 4548
rect 16114 4536 16120 4548
rect 13688 4508 16120 4536
rect 13688 4496 13694 4508
rect 16114 4496 16120 4508
rect 16172 4496 16178 4548
rect 16224 4536 16252 4576
rect 17221 4573 17233 4607
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18138 4604 18144 4616
rect 18095 4576 18144 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 17865 4539 17923 4545
rect 17865 4536 17877 4539
rect 16224 4508 17877 4536
rect 17865 4505 17877 4508
rect 17911 4505 17923 4539
rect 17865 4499 17923 4505
rect 4430 4428 4436 4480
rect 4488 4428 4494 4480
rect 5077 4471 5135 4477
rect 5077 4437 5089 4471
rect 5123 4468 5135 4471
rect 5258 4468 5264 4480
rect 5123 4440 5264 4468
rect 5123 4437 5135 4440
rect 5077 4431 5135 4437
rect 5258 4428 5264 4440
rect 5316 4468 5322 4480
rect 5629 4471 5687 4477
rect 5629 4468 5641 4471
rect 5316 4440 5641 4468
rect 5316 4428 5322 4440
rect 5629 4437 5641 4440
rect 5675 4437 5687 4471
rect 5629 4431 5687 4437
rect 7996 4471 8054 4477
rect 7996 4437 8008 4471
rect 8042 4468 8054 4471
rect 17494 4468 17500 4480
rect 8042 4440 17500 4468
rect 8042 4437 8054 4440
rect 7996 4431 8054 4437
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 1104 4378 18860 4400
rect 1104 4326 3829 4378
rect 3881 4326 3893 4378
rect 3945 4326 3957 4378
rect 4009 4326 4021 4378
rect 4073 4326 4085 4378
rect 4137 4326 8268 4378
rect 8320 4326 8332 4378
rect 8384 4326 8396 4378
rect 8448 4326 8460 4378
rect 8512 4326 8524 4378
rect 8576 4326 12707 4378
rect 12759 4326 12771 4378
rect 12823 4326 12835 4378
rect 12887 4326 12899 4378
rect 12951 4326 12963 4378
rect 13015 4326 17146 4378
rect 17198 4326 17210 4378
rect 17262 4326 17274 4378
rect 17326 4326 17338 4378
rect 17390 4326 17402 4378
rect 17454 4326 18860 4378
rect 1104 4304 18860 4326
rect 1854 4224 1860 4276
rect 1912 4264 1918 4276
rect 1949 4267 2007 4273
rect 1949 4264 1961 4267
rect 1912 4236 1961 4264
rect 1912 4224 1918 4236
rect 1949 4233 1961 4236
rect 1995 4264 2007 4267
rect 3326 4264 3332 4276
rect 1995 4236 3332 4264
rect 1995 4233 2007 4236
rect 1949 4227 2007 4233
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 4338 4264 4344 4276
rect 4172 4236 4344 4264
rect 4172 4196 4200 4236
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 8846 4264 8852 4276
rect 4488 4236 8852 4264
rect 4488 4224 4494 4236
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 9824 4236 11008 4264
rect 9824 4224 9830 4236
rect 5353 4199 5411 4205
rect 4094 4168 4200 4196
rect 4816 4168 5028 4196
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 2700 4060 2728 4091
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2832 4100 2973 4128
rect 2832 4088 2838 4100
rect 2961 4097 2973 4100
rect 3007 4097 3019 4131
rect 4816 4128 4844 4168
rect 2961 4091 3019 4097
rect 4356 4100 4844 4128
rect 4356 4060 4384 4100
rect 4890 4088 4896 4140
rect 4948 4088 4954 4140
rect 5000 4128 5028 4168
rect 5353 4165 5365 4199
rect 5399 4196 5411 4199
rect 5534 4196 5540 4208
rect 5399 4168 5540 4196
rect 5399 4165 5411 4168
rect 5353 4159 5411 4165
rect 5534 4156 5540 4168
rect 5592 4156 5598 4208
rect 10778 4196 10784 4208
rect 10350 4168 10784 4196
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 10980 4196 11008 4236
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 13872 4236 14320 4264
rect 13872 4224 13878 4236
rect 14292 4196 14320 4236
rect 15102 4196 15108 4208
rect 10980 4168 11100 4196
rect 14214 4168 15108 4196
rect 5721 4131 5779 4137
rect 5000 4100 5488 4128
rect 2547 4032 4384 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 4430 4020 4436 4072
rect 4488 4020 4494 4072
rect 4795 4063 4853 4069
rect 4795 4029 4807 4063
rect 4841 4029 4853 4063
rect 5460 4060 5488 4100
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 5767 4100 6193 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 6181 4097 6193 4100
rect 6227 4128 6239 4131
rect 6270 4128 6276 4140
rect 6227 4100 6276 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 8938 4128 8944 4140
rect 7524 4100 8944 4128
rect 7524 4088 7530 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 11072 4137 11100 4168
rect 15102 4156 15108 4168
rect 15160 4156 15166 4208
rect 17402 4156 17408 4208
rect 17460 4156 17466 4208
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4128 11115 4131
rect 13078 4128 13084 4140
rect 11103 4100 13084 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 13078 4088 13084 4100
rect 13136 4128 13142 4140
rect 13136 4100 13492 4128
rect 13136 4088 13142 4100
rect 10781 4063 10839 4069
rect 5460 4032 9444 4060
rect 4795 4023 4853 4029
rect 750 3952 756 4004
rect 808 3992 814 4004
rect 2869 3995 2927 4001
rect 2869 3992 2881 3995
rect 808 3964 2881 3992
rect 808 3952 814 3964
rect 2869 3961 2881 3964
rect 2915 3961 2927 3995
rect 2869 3955 2927 3961
rect 4816 3992 4844 4023
rect 6178 3992 6184 4004
rect 4816 3964 6184 3992
rect 3510 3884 3516 3936
rect 3568 3924 3574 3936
rect 4816 3924 4844 3964
rect 6178 3952 6184 3964
rect 6236 3952 6242 4004
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 9088 3964 9321 3992
rect 9088 3952 9094 3964
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 3568 3896 4844 3924
rect 9416 3924 9444 4032
rect 10781 4029 10793 4063
rect 10827 4060 10839 4063
rect 12618 4060 12624 4072
rect 10827 4032 12624 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 12894 4020 12900 4072
rect 12952 4020 12958 4072
rect 11146 3924 11152 3936
rect 9416 3896 11152 3924
rect 3568 3884 3574 3896
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 11664 3896 12817 3924
rect 11664 3884 11670 3896
rect 12805 3893 12817 3896
rect 12851 3924 12863 3927
rect 13354 3924 13360 3936
rect 12851 3896 13360 3924
rect 12851 3893 12863 3896
rect 12805 3887 12863 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 13464 3924 13492 4100
rect 15286 4088 15292 4140
rect 15344 4088 15350 4140
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 15565 4131 15623 4137
rect 15565 4128 15577 4131
rect 15528 4100 15577 4128
rect 15528 4088 15534 4100
rect 15565 4097 15577 4100
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 17037 4131 17095 4137
rect 17037 4128 17049 4131
rect 16448 4100 17049 4128
rect 16448 4088 16454 4100
rect 17037 4097 17049 4100
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 17920 4100 18521 4128
rect 17920 4088 17926 4100
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 14332 4032 14657 4060
rect 14332 4020 14338 4032
rect 14645 4029 14657 4032
rect 14691 4029 14703 4063
rect 14645 4023 14703 4029
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4060 14979 4063
rect 16298 4060 16304 4072
rect 14967 4032 16304 4060
rect 14967 4029 14979 4032
rect 14921 4023 14979 4029
rect 14936 3924 14964 4023
rect 16298 4020 16304 4032
rect 16356 4060 16362 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16356 4032 16681 4060
rect 16356 4020 16362 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 13464 3896 14964 3924
rect 16390 3884 16396 3936
rect 16448 3884 16454 3936
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3016 3692 4384 3720
rect 3016 3680 3022 3692
rect 2685 3655 2743 3661
rect 2685 3621 2697 3655
rect 2731 3652 2743 3655
rect 3694 3652 3700 3664
rect 2731 3624 3700 3652
rect 2731 3621 2743 3624
rect 2685 3615 2743 3621
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 4356 3652 4384 3692
rect 4430 3680 4436 3732
rect 4488 3720 4494 3732
rect 4893 3723 4951 3729
rect 4893 3720 4905 3723
rect 4488 3692 4905 3720
rect 4488 3680 4494 3692
rect 4893 3689 4905 3692
rect 4939 3689 4951 3723
rect 4893 3683 4951 3689
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 6454 3720 6460 3732
rect 5776 3692 6460 3720
rect 5776 3680 5782 3692
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 9861 3723 9919 3729
rect 9861 3720 9873 3723
rect 8128 3692 9873 3720
rect 8128 3652 8156 3692
rect 9861 3689 9873 3692
rect 9907 3720 9919 3723
rect 10042 3720 10048 3732
rect 9907 3692 10048 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10410 3680 10416 3732
rect 10468 3720 10474 3732
rect 11146 3720 11152 3732
rect 10468 3692 11152 3720
rect 10468 3680 10474 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 11388 3692 12848 3720
rect 11388 3680 11394 3692
rect 4356 3624 8156 3652
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 9585 3655 9643 3661
rect 9585 3652 9597 3655
rect 8812 3624 9597 3652
rect 8812 3612 8818 3624
rect 9585 3621 9597 3624
rect 9631 3652 9643 3655
rect 12342 3652 12348 3664
rect 9631 3624 12348 3652
rect 9631 3621 9643 3624
rect 9585 3615 9643 3621
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 842 3544 848 3596
rect 900 3584 906 3596
rect 1581 3587 1639 3593
rect 1581 3584 1593 3587
rect 900 3556 1593 3584
rect 900 3544 906 3556
rect 1581 3553 1593 3556
rect 1627 3553 1639 3587
rect 2958 3584 2964 3596
rect 1581 3547 1639 3553
rect 1872 3556 2964 3584
rect 1872 3525 1900 3556
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 3605 3587 3663 3593
rect 3605 3553 3617 3587
rect 3651 3584 3663 3587
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 3651 3556 4169 3584
rect 3651 3553 3663 3556
rect 3605 3547 3663 3553
rect 4157 3553 4169 3556
rect 4203 3584 4215 3587
rect 11790 3584 11796 3596
rect 4203 3556 11796 3584
rect 4203 3553 4215 3556
rect 4157 3547 4215 3553
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 12820 3593 12848 3692
rect 13630 3680 13636 3732
rect 13688 3680 13694 3732
rect 15010 3720 15016 3732
rect 13740 3692 15016 3720
rect 13170 3612 13176 3664
rect 13228 3652 13234 3664
rect 13740 3652 13768 3692
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 15194 3680 15200 3732
rect 15252 3680 15258 3732
rect 15470 3680 15476 3732
rect 15528 3680 15534 3732
rect 13228 3624 13768 3652
rect 13228 3612 13234 3624
rect 14642 3612 14648 3664
rect 14700 3612 14706 3664
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 12851 3556 13308 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 3050 3516 3056 3528
rect 2547 3488 3056 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4525 3519 4583 3525
rect 4525 3485 4537 3519
rect 4571 3516 4583 3519
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 4571 3488 5365 3516
rect 4571 3485 4583 3488
rect 4525 3479 4583 3485
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 5353 3479 5411 3485
rect 4356 3448 4384 3479
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 5920 3448 5948 3479
rect 8018 3476 8024 3528
rect 8076 3476 8082 3528
rect 8662 3476 8668 3528
rect 8720 3476 8726 3528
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 12618 3516 12624 3528
rect 10744 3488 12624 3516
rect 10744 3476 10750 3488
rect 12618 3476 12624 3488
rect 12676 3516 12682 3528
rect 13280 3525 13308 3556
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 13412 3556 13497 3584
rect 13412 3544 13418 3556
rect 13469 3525 13497 3556
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 14277 3587 14335 3593
rect 14277 3584 14289 3587
rect 13780 3556 14289 3584
rect 13780 3544 13786 3556
rect 14277 3553 14289 3556
rect 14323 3584 14335 3587
rect 14458 3584 14464 3596
rect 14323 3556 14464 3584
rect 14323 3553 14335 3556
rect 14277 3547 14335 3553
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 14921 3587 14979 3593
rect 14921 3553 14933 3587
rect 14967 3584 14979 3587
rect 15212 3584 15240 3680
rect 14967 3556 15240 3584
rect 14967 3553 14979 3556
rect 14921 3547 14979 3553
rect 15838 3544 15844 3596
rect 15896 3584 15902 3596
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15896 3556 16037 3584
rect 15896 3544 15902 3556
rect 16025 3553 16037 3556
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 16298 3544 16304 3596
rect 16356 3544 16362 3596
rect 18046 3544 18052 3596
rect 18104 3544 18110 3596
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 12676 3488 13093 3516
rect 12676 3476 12682 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13265 3519 13323 3525
rect 13265 3485 13277 3519
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 13454 3519 13512 3525
rect 13454 3485 13466 3519
rect 13500 3485 13512 3519
rect 13454 3479 13512 3485
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 4356 3420 4568 3448
rect 4540 3392 4568 3420
rect 5368 3420 5948 3448
rect 5368 3392 5396 3420
rect 6086 3408 6092 3460
rect 6144 3408 6150 3460
rect 6270 3408 6276 3460
rect 6328 3448 6334 3460
rect 8680 3448 8708 3476
rect 6328 3420 8708 3448
rect 6328 3408 6334 3420
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 10778 3448 10784 3460
rect 10100 3420 10784 3448
rect 10100 3408 10106 3420
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 13357 3451 13415 3457
rect 11204 3420 13216 3448
rect 11204 3408 11210 3420
rect 2130 3340 2136 3392
rect 2188 3340 2194 3392
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 3973 3383 4031 3389
rect 3973 3380 3985 3383
rect 2556 3352 3985 3380
rect 2556 3340 2562 3352
rect 3973 3349 3985 3352
rect 4019 3380 4031 3383
rect 4430 3380 4436 3392
rect 4019 3352 4436 3380
rect 4019 3349 4031 3352
rect 3973 3343 4031 3349
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 4522 3340 4528 3392
rect 4580 3340 4586 3392
rect 5350 3340 5356 3392
rect 5408 3340 5414 3392
rect 7834 3340 7840 3392
rect 7892 3340 7898 3392
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8662 3380 8668 3392
rect 8527 3352 8668 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 9030 3340 9036 3392
rect 9088 3380 9094 3392
rect 9125 3383 9183 3389
rect 9125 3380 9137 3383
rect 9088 3352 9137 3380
rect 9088 3340 9094 3352
rect 9125 3349 9137 3352
rect 9171 3349 9183 3383
rect 9125 3343 9183 3349
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 12342 3380 12348 3392
rect 12299 3352 12348 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 13188 3380 13216 3420
rect 13357 3417 13369 3451
rect 13403 3448 13415 3451
rect 14090 3448 14096 3460
rect 13403 3420 14096 3448
rect 13403 3417 13415 3420
rect 13357 3411 13415 3417
rect 14090 3408 14096 3420
rect 14148 3408 14154 3460
rect 14384 3380 14412 3479
rect 16206 3476 16212 3528
rect 16264 3516 16270 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16264 3488 16681 3516
rect 16264 3476 16270 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 15841 3451 15899 3457
rect 15841 3448 15853 3451
rect 15620 3420 15853 3448
rect 15620 3408 15626 3420
rect 15841 3417 15853 3420
rect 15887 3417 15899 3451
rect 15841 3411 15899 3417
rect 16960 3420 17066 3448
rect 13188 3352 14412 3380
rect 15930 3340 15936 3392
rect 15988 3340 15994 3392
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 16960 3380 16988 3420
rect 17402 3380 17408 3392
rect 16448 3352 17408 3380
rect 16448 3340 16454 3352
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 1104 3290 18860 3312
rect 1104 3238 3829 3290
rect 3881 3238 3893 3290
rect 3945 3238 3957 3290
rect 4009 3238 4021 3290
rect 4073 3238 4085 3290
rect 4137 3238 8268 3290
rect 8320 3238 8332 3290
rect 8384 3238 8396 3290
rect 8448 3238 8460 3290
rect 8512 3238 8524 3290
rect 8576 3238 12707 3290
rect 12759 3238 12771 3290
rect 12823 3238 12835 3290
rect 12887 3238 12899 3290
rect 12951 3238 12963 3290
rect 13015 3238 17146 3290
rect 17198 3238 17210 3290
rect 17262 3238 17274 3290
rect 17326 3238 17338 3290
rect 17390 3238 17402 3290
rect 17454 3238 18860 3290
rect 1104 3216 18860 3238
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 1949 3179 2007 3185
rect 1949 3176 1961 3179
rect 1820 3148 1961 3176
rect 1820 3136 1826 3148
rect 1949 3145 1961 3148
rect 1995 3145 2007 3179
rect 1949 3139 2007 3145
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3602 3176 3608 3188
rect 3200 3148 3608 3176
rect 3200 3136 3206 3148
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 4249 3179 4307 3185
rect 4249 3145 4261 3179
rect 4295 3176 4307 3179
rect 4522 3176 4528 3188
rect 4295 3148 4528 3176
rect 4295 3145 4307 3148
rect 4249 3139 4307 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 4890 3176 4896 3188
rect 4663 3148 4896 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 5261 3179 5319 3185
rect 5261 3145 5273 3179
rect 5307 3176 5319 3179
rect 5350 3176 5356 3188
rect 5307 3148 5356 3176
rect 5307 3145 5319 3148
rect 5261 3139 5319 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5592 3148 5641 3176
rect 5592 3136 5598 3148
rect 5629 3145 5641 3148
rect 5675 3176 5687 3179
rect 5994 3176 6000 3188
rect 5675 3148 6000 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 7466 3136 7472 3188
rect 7524 3136 7530 3188
rect 10134 3136 10140 3188
rect 10192 3136 10198 3188
rect 10318 3136 10324 3188
rect 10376 3136 10382 3188
rect 12526 3136 12532 3188
rect 12584 3136 12590 3188
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 13354 3176 13360 3188
rect 12676 3148 13360 3176
rect 12676 3136 12682 3148
rect 13354 3136 13360 3148
rect 13412 3176 13418 3188
rect 15286 3176 15292 3188
rect 13412 3148 15292 3176
rect 13412 3136 13418 3148
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15838 3136 15844 3188
rect 15896 3176 15902 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 15896 3148 16865 3176
rect 15896 3136 15902 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 17770 3136 17776 3188
rect 17828 3136 17834 3188
rect 1872 3080 3556 3108
rect 1872 3049 1900 3080
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2130 3000 2136 3052
rect 2188 3000 2194 3052
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2682 3040 2688 3052
rect 2639 3012 2688 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 2823 3012 3464 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 842 2932 848 2984
rect 900 2972 906 2984
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 900 2944 1593 2972
rect 900 2932 906 2944
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 2700 2972 2728 3000
rect 3053 2975 3111 2981
rect 3053 2972 3065 2975
rect 2700 2944 3065 2972
rect 1581 2935 1639 2941
rect 3053 2941 3065 2944
rect 3099 2941 3111 2975
rect 3053 2935 3111 2941
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2904 2467 2907
rect 3142 2904 3148 2916
rect 2455 2876 3148 2904
rect 2455 2873 2467 2876
rect 2409 2867 2467 2873
rect 3142 2864 3148 2876
rect 3200 2864 3206 2916
rect 3436 2904 3464 3012
rect 3528 2981 3556 3080
rect 7926 3068 7932 3120
rect 7984 3108 7990 3120
rect 14918 3108 14924 3120
rect 7984 3080 10640 3108
rect 14306 3080 14924 3108
rect 7984 3068 7990 3080
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 5500 3012 7849 3040
rect 5500 3000 5506 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 6270 2972 6276 2984
rect 3559 2944 6276 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 7374 2932 7380 2984
rect 7432 2972 7438 2984
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7432 2944 7573 2972
rect 7432 2932 7438 2944
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 7852 2972 7880 3003
rect 8110 3000 8116 3052
rect 8168 3000 8174 3052
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3040 8723 3043
rect 8754 3040 8760 3052
rect 8711 3012 8760 3040
rect 8711 3009 8723 3012
rect 8665 3003 8723 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 8938 3000 8944 3052
rect 8996 3000 9002 3052
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 10612 3049 10640 3080
rect 14918 3068 14924 3080
rect 14976 3108 14982 3120
rect 15657 3111 15715 3117
rect 15657 3108 15669 3111
rect 14976 3080 15669 3108
rect 14976 3068 14982 3080
rect 15657 3077 15669 3080
rect 15703 3108 15715 3111
rect 16117 3111 16175 3117
rect 16117 3108 16129 3111
rect 15703 3080 16129 3108
rect 15703 3077 15715 3080
rect 15657 3071 15715 3077
rect 16117 3077 16129 3080
rect 16163 3108 16175 3111
rect 16390 3108 16396 3120
rect 16163 3080 16396 3108
rect 16163 3077 16175 3080
rect 16117 3071 16175 3077
rect 16390 3068 16396 3080
rect 16448 3068 16454 3120
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 9640 3012 10517 3040
rect 9640 3000 9646 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 10686 3000 10692 3052
rect 10744 3000 10750 3052
rect 10778 3000 10784 3052
rect 10836 3000 10842 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10888 3012 10977 3040
rect 8294 2972 8300 2984
rect 7852 2944 8300 2972
rect 7561 2935 7619 2941
rect 8294 2932 8300 2944
rect 8352 2932 8358 2984
rect 9401 2975 9459 2981
rect 9401 2941 9413 2975
rect 9447 2972 9459 2975
rect 9674 2972 9680 2984
rect 9447 2944 9680 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 10318 2972 10324 2984
rect 9815 2944 10324 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 9858 2904 9864 2916
rect 3436 2876 9864 2904
rect 9858 2864 9864 2876
rect 9916 2864 9922 2916
rect 10134 2864 10140 2916
rect 10192 2904 10198 2916
rect 10888 2904 10916 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 11606 2932 11612 2984
rect 11664 2972 11670 2984
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11664 2944 11897 2972
rect 11664 2932 11670 2944
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 12176 2972 12204 3003
rect 12342 3000 12348 3052
rect 12400 3000 12406 3052
rect 13170 3040 13176 3052
rect 12452 3012 13176 3040
rect 12452 2972 12480 3012
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3040 17371 3043
rect 18233 3043 18291 3049
rect 17359 3012 18184 3040
rect 17359 3009 17371 3012
rect 17313 3003 17371 3009
rect 12176 2944 12480 2972
rect 11885 2935 11943 2941
rect 12618 2932 12624 2984
rect 12676 2972 12682 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12676 2944 12909 2972
rect 12676 2932 12682 2944
rect 12897 2941 12909 2944
rect 12943 2972 12955 2975
rect 13078 2972 13084 2984
rect 12943 2944 13084 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13265 2975 13323 2981
rect 13265 2941 13277 2975
rect 13311 2972 13323 2975
rect 13446 2972 13452 2984
rect 13311 2944 13452 2972
rect 13311 2941 13323 2944
rect 13265 2935 13323 2941
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 14090 2932 14096 2984
rect 14148 2972 14154 2984
rect 14645 2975 14703 2981
rect 14645 2972 14657 2975
rect 14148 2944 14657 2972
rect 14148 2932 14154 2944
rect 14645 2941 14657 2944
rect 14691 2941 14703 2975
rect 14645 2935 14703 2941
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 18156 2981 18184 3012
rect 18233 3009 18245 3043
rect 18279 3040 18291 3043
rect 18414 3040 18420 3052
rect 18279 3012 18420 3040
rect 18279 3009 18291 3012
rect 18233 3003 18291 3009
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 17957 2975 18015 2981
rect 17957 2972 17969 2975
rect 17460 2944 17969 2972
rect 17460 2932 17466 2944
rect 17957 2941 17969 2944
rect 18003 2941 18015 2975
rect 17957 2935 18015 2941
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2972 18199 2975
rect 19334 2972 19340 2984
rect 18187 2944 19340 2972
rect 18187 2941 18199 2944
rect 18141 2935 18199 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 15930 2904 15936 2916
rect 10192 2876 10916 2904
rect 10980 2876 12940 2904
rect 10192 2864 10198 2876
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 8754 2836 8760 2848
rect 6880 2808 8760 2836
rect 6880 2796 6886 2808
rect 8754 2796 8760 2808
rect 8812 2836 8818 2848
rect 10980 2836 11008 2876
rect 8812 2808 11008 2836
rect 8812 2796 8818 2808
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11241 2839 11299 2845
rect 11241 2836 11253 2839
rect 11112 2808 11253 2836
rect 11112 2796 11118 2808
rect 11241 2805 11253 2808
rect 11287 2805 11299 2839
rect 12912 2836 12940 2876
rect 15304 2876 15936 2904
rect 15304 2845 15332 2876
rect 15930 2864 15936 2876
rect 15988 2864 15994 2916
rect 15289 2839 15347 2845
rect 15289 2836 15301 2839
rect 12912 2808 15301 2836
rect 11241 2799 11299 2805
rect 15289 2805 15301 2808
rect 15335 2805 15347 2839
rect 15289 2799 15347 2805
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 1486 2592 1492 2644
rect 1544 2632 1550 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 1544 2604 2421 2632
rect 1544 2592 1550 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2409 2595 2467 2601
rect 4430 2592 4436 2644
rect 4488 2592 4494 2644
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 7285 2635 7343 2641
rect 7285 2632 7297 2635
rect 6604 2604 7297 2632
rect 6604 2592 6610 2604
rect 7285 2601 7297 2604
rect 7331 2601 7343 2635
rect 7285 2595 7343 2601
rect 934 2524 940 2576
rect 992 2564 998 2576
rect 2133 2567 2191 2573
rect 2133 2564 2145 2567
rect 992 2536 2145 2564
rect 992 2524 998 2536
rect 2133 2533 2145 2536
rect 2179 2533 2191 2567
rect 7190 2564 7196 2576
rect 2133 2527 2191 2533
rect 6104 2536 7196 2564
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 4111 2468 5917 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 5905 2465 5917 2468
rect 5951 2496 5963 2499
rect 6104 2496 6132 2536
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 5951 2468 6132 2496
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 7300 2496 7328 2595
rect 7466 2592 7472 2644
rect 7524 2592 7530 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 10226 2632 10232 2644
rect 8527 2604 10232 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10594 2592 10600 2644
rect 10652 2592 10658 2644
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 11146 2632 11152 2644
rect 11103 2604 11152 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11900 2604 13308 2632
rect 7484 2564 7512 2592
rect 7484 2536 8064 2564
rect 8036 2505 8064 2536
rect 8754 2524 8760 2576
rect 8812 2524 8818 2576
rect 8938 2524 8944 2576
rect 8996 2564 9002 2576
rect 11900 2564 11928 2604
rect 8996 2536 11928 2564
rect 13280 2564 13308 2604
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13541 2635 13599 2641
rect 13541 2632 13553 2635
rect 13412 2604 13553 2632
rect 13412 2592 13418 2604
rect 13541 2601 13553 2604
rect 13587 2601 13599 2635
rect 13998 2632 14004 2644
rect 13541 2595 13599 2601
rect 13648 2604 14004 2632
rect 13648 2564 13676 2604
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 14424 2604 14964 2632
rect 14424 2592 14430 2604
rect 14936 2576 14964 2604
rect 17310 2592 17316 2644
rect 17368 2592 17374 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 18598 2632 18604 2644
rect 17819 2604 18604 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 13280 2536 13676 2564
rect 8996 2524 9002 2536
rect 14458 2524 14464 2576
rect 14516 2564 14522 2576
rect 14553 2567 14611 2573
rect 14553 2564 14565 2567
rect 14516 2536 14565 2564
rect 14516 2524 14522 2536
rect 14553 2533 14565 2536
rect 14599 2533 14611 2567
rect 14553 2527 14611 2533
rect 14918 2524 14924 2576
rect 14976 2564 14982 2576
rect 15381 2567 15439 2573
rect 14976 2536 15332 2564
rect 14976 2524 14982 2536
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7300 2468 7849 2496
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2465 8079 2499
rect 8021 2459 8079 2465
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 11793 2499 11851 2505
rect 8352 2468 10088 2496
rect 8352 2456 8358 2468
rect 1854 2388 1860 2440
rect 1912 2388 1918 2440
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2866 2428 2872 2440
rect 2639 2400 2872 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 842 2320 848 2372
rect 900 2360 906 2372
rect 1581 2363 1639 2369
rect 1581 2360 1593 2363
rect 900 2332 1593 2360
rect 900 2320 906 2332
rect 1581 2329 1593 2332
rect 1627 2329 1639 2363
rect 1964 2360 1992 2391
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 6687 2400 7665 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 7653 2397 7665 2400
rect 7699 2428 7711 2431
rect 7742 2428 7748 2440
rect 7699 2400 7748 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8662 2428 8668 2440
rect 8619 2400 8668 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 2774 2360 2780 2372
rect 1964 2332 2780 2360
rect 1581 2323 1639 2329
rect 2774 2320 2780 2332
rect 2832 2360 2838 2372
rect 3237 2363 3295 2369
rect 3237 2360 3249 2363
rect 2832 2332 3249 2360
rect 2832 2320 2838 2332
rect 3237 2329 3249 2332
rect 3283 2329 3295 2363
rect 3237 2323 3295 2329
rect 6886 2332 9352 2360
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 6886 2292 6914 2332
rect 5316 2264 6914 2292
rect 7009 2295 7067 2301
rect 5316 2252 5322 2264
rect 7009 2261 7021 2295
rect 7055 2292 7067 2295
rect 8113 2295 8171 2301
rect 8113 2292 8125 2295
rect 7055 2264 8125 2292
rect 7055 2261 7067 2264
rect 7009 2255 7067 2261
rect 8113 2261 8125 2264
rect 8159 2292 8171 2295
rect 9214 2292 9220 2304
rect 8159 2264 9220 2292
rect 8159 2261 8171 2264
rect 8113 2255 8171 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9324 2301 9352 2332
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 9950 2252 9956 2304
rect 10008 2252 10014 2304
rect 10060 2292 10088 2468
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 12618 2496 12624 2508
rect 11839 2468 12624 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 12860 2468 15240 2496
rect 12860 2456 12866 2468
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10376 2400 10425 2428
rect 10376 2388 10382 2400
rect 10413 2397 10425 2400
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11112 2400 11253 2428
rect 11112 2388 11118 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 12066 2320 12072 2372
rect 12124 2320 12130 2372
rect 13814 2360 13820 2372
rect 13294 2332 13820 2360
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 12802 2292 12808 2304
rect 10060 2264 12808 2292
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 13354 2252 13360 2304
rect 13412 2292 13418 2304
rect 14093 2295 14151 2301
rect 14093 2292 14105 2295
rect 13412 2264 14105 2292
rect 13412 2252 13418 2264
rect 14093 2261 14105 2264
rect 14139 2261 14151 2295
rect 14292 2292 14320 2391
rect 14550 2388 14556 2440
rect 14608 2428 14614 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14608 2400 14841 2428
rect 14608 2388 14614 2400
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 14844 2360 14872 2391
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 15102 2388 15108 2440
rect 15160 2388 15166 2440
rect 15212 2437 15240 2468
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 15304 2428 15332 2536
rect 15381 2533 15393 2567
rect 15427 2564 15439 2567
rect 18230 2564 18236 2576
rect 15427 2536 18236 2564
rect 15427 2533 15439 2536
rect 15381 2527 15439 2533
rect 18230 2524 18236 2536
rect 18288 2524 18294 2576
rect 19426 2428 19432 2440
rect 15304 2400 19432 2428
rect 15197 2391 15255 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 14844 2332 15761 2360
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 18782 2360 18788 2372
rect 15749 2323 15807 2329
rect 17236 2332 18788 2360
rect 17236 2292 17264 2332
rect 18782 2320 18788 2332
rect 18840 2320 18846 2372
rect 14292 2264 17264 2292
rect 14093 2255 14151 2261
rect 1104 2202 18860 2224
rect 1104 2150 3829 2202
rect 3881 2150 3893 2202
rect 3945 2150 3957 2202
rect 4009 2150 4021 2202
rect 4073 2150 4085 2202
rect 4137 2150 8268 2202
rect 8320 2150 8332 2202
rect 8384 2150 8396 2202
rect 8448 2150 8460 2202
rect 8512 2150 8524 2202
rect 8576 2150 12707 2202
rect 12759 2150 12771 2202
rect 12823 2150 12835 2202
rect 12887 2150 12899 2202
rect 12951 2150 12963 2202
rect 13015 2150 17146 2202
rect 17198 2150 17210 2202
rect 17262 2150 17274 2202
rect 17326 2150 17338 2202
rect 17390 2150 17402 2202
rect 17454 2150 18860 2202
rect 1104 2128 18860 2150
rect 8110 2048 8116 2100
rect 8168 2088 8174 2100
rect 15102 2088 15108 2100
rect 8168 2060 15108 2088
rect 8168 2048 8174 2060
rect 15102 2048 15108 2060
rect 15160 2048 15166 2100
rect 9214 1980 9220 2032
rect 9272 2020 9278 2032
rect 11698 2020 11704 2032
rect 9272 1992 11704 2020
rect 9272 1980 9278 1992
rect 11698 1980 11704 1992
rect 11756 1980 11762 2032
rect 7190 1912 7196 1964
rect 7248 1952 7254 1964
rect 11238 1952 11244 1964
rect 7248 1924 11244 1952
rect 7248 1912 7254 1924
rect 11238 1912 11244 1924
rect 11296 1912 11302 1964
rect 566 1844 572 1896
rect 624 1884 630 1896
rect 12066 1884 12072 1896
rect 624 1856 12072 1884
rect 624 1844 630 1856
rect 12066 1844 12072 1856
rect 12124 1844 12130 1896
<< via1 >>
rect 6184 17620 6236 17672
rect 13820 17620 13872 17672
rect 7380 17552 7432 17604
rect 18972 17552 19024 17604
rect 6000 17484 6052 17536
rect 13084 17484 13136 17536
rect 3829 17382 3881 17434
rect 3893 17382 3945 17434
rect 3957 17382 4009 17434
rect 4021 17382 4073 17434
rect 4085 17382 4137 17434
rect 8268 17382 8320 17434
rect 8332 17382 8384 17434
rect 8396 17382 8448 17434
rect 8460 17382 8512 17434
rect 8524 17382 8576 17434
rect 12707 17382 12759 17434
rect 12771 17382 12823 17434
rect 12835 17382 12887 17434
rect 12899 17382 12951 17434
rect 12963 17382 13015 17434
rect 17146 17382 17198 17434
rect 17210 17382 17262 17434
rect 17274 17382 17326 17434
rect 17338 17382 17390 17434
rect 17402 17382 17454 17434
rect 3700 17280 3752 17332
rect 1492 17144 1544 17196
rect 2872 17212 2924 17264
rect 2964 17212 3016 17264
rect 3608 17212 3660 17264
rect 4344 17212 4396 17264
rect 6828 17280 6880 17332
rect 7380 17323 7432 17332
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6552 17187 6604 17196
rect 6552 17153 6601 17187
rect 6601 17153 6604 17187
rect 6552 17144 6604 17153
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 9220 17280 9272 17332
rect 7564 17212 7616 17264
rect 16948 17280 17000 17332
rect 9404 17212 9456 17264
rect 2688 17076 2740 17128
rect 3516 17076 3568 17128
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 5632 17119 5684 17128
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 7196 17144 7248 17196
rect 7656 17144 7708 17196
rect 9772 17144 9824 17196
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 12164 17255 12216 17264
rect 12164 17221 12173 17255
rect 12173 17221 12207 17255
rect 12207 17221 12216 17255
rect 12164 17212 12216 17221
rect 12532 17212 12584 17264
rect 15200 17212 15252 17264
rect 13636 17144 13688 17196
rect 8392 17076 8444 17128
rect 8760 17076 8812 17128
rect 16028 17076 16080 17128
rect 1952 17008 2004 17060
rect 2688 16940 2740 16992
rect 3056 16940 3108 16992
rect 3792 16940 3844 16992
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 6000 17008 6052 17060
rect 11152 17008 11204 17060
rect 5908 16940 5960 16992
rect 6552 16940 6604 16992
rect 7104 16940 7156 16992
rect 7380 16940 7432 16992
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 8852 16940 8904 16992
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9128 16940 9180 16949
rect 10784 16940 10836 16992
rect 11796 16940 11848 16992
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 13636 16940 13688 16992
rect 16304 16983 16356 16992
rect 16304 16949 16313 16983
rect 16313 16949 16347 16983
rect 16347 16949 16356 16983
rect 16304 16940 16356 16949
rect 3169 16838 3221 16890
rect 3233 16838 3285 16890
rect 3297 16838 3349 16890
rect 3361 16838 3413 16890
rect 3425 16838 3477 16890
rect 7608 16838 7660 16890
rect 7672 16838 7724 16890
rect 7736 16838 7788 16890
rect 7800 16838 7852 16890
rect 7864 16838 7916 16890
rect 12047 16838 12099 16890
rect 12111 16838 12163 16890
rect 12175 16838 12227 16890
rect 12239 16838 12291 16890
rect 12303 16838 12355 16890
rect 16486 16838 16538 16890
rect 16550 16838 16602 16890
rect 16614 16838 16666 16890
rect 16678 16838 16730 16890
rect 16742 16838 16794 16890
rect 4436 16736 4488 16788
rect 2044 16643 2096 16652
rect 2044 16609 2053 16643
rect 2053 16609 2087 16643
rect 2087 16609 2096 16643
rect 2044 16600 2096 16609
rect 1952 16532 2004 16584
rect 2964 16600 3016 16652
rect 3792 16668 3844 16720
rect 4344 16668 4396 16720
rect 5540 16736 5592 16788
rect 5816 16779 5868 16788
rect 5816 16745 5825 16779
rect 5825 16745 5859 16779
rect 5859 16745 5868 16779
rect 5816 16736 5868 16745
rect 6000 16736 6052 16788
rect 6920 16736 6972 16788
rect 7288 16779 7340 16788
rect 7288 16745 7297 16779
rect 7297 16745 7331 16779
rect 7331 16745 7340 16779
rect 7288 16736 7340 16745
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 2780 16532 2832 16584
rect 4252 16600 4304 16652
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 5540 16600 5592 16652
rect 8484 16600 8536 16652
rect 8944 16600 8996 16652
rect 11244 16736 11296 16788
rect 12072 16736 12124 16788
rect 9496 16668 9548 16720
rect 11520 16668 11572 16720
rect 12256 16668 12308 16720
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 16304 16736 16356 16788
rect 9128 16600 9180 16652
rect 6644 16532 6696 16584
rect 8668 16532 8720 16584
rect 2228 16464 2280 16516
rect 1860 16396 1912 16448
rect 2780 16396 2832 16448
rect 4620 16439 4672 16448
rect 4620 16405 4629 16439
rect 4629 16405 4663 16439
rect 4663 16405 4672 16439
rect 4620 16396 4672 16405
rect 5264 16464 5316 16516
rect 8484 16464 8536 16516
rect 9312 16575 9364 16584
rect 9312 16541 9321 16575
rect 9321 16541 9355 16575
rect 9355 16541 9364 16575
rect 9312 16532 9364 16541
rect 13820 16711 13872 16720
rect 13820 16677 13829 16711
rect 13829 16677 13863 16711
rect 13863 16677 13872 16711
rect 13820 16668 13872 16677
rect 9680 16532 9732 16584
rect 10140 16532 10192 16584
rect 5448 16396 5500 16448
rect 6644 16396 6696 16448
rect 9128 16396 9180 16448
rect 11060 16464 11112 16516
rect 11980 16532 12032 16584
rect 12072 16575 12124 16584
rect 12072 16541 12081 16575
rect 12081 16541 12115 16575
rect 12115 16541 12124 16575
rect 12072 16532 12124 16541
rect 14740 16600 14792 16652
rect 15200 16600 15252 16652
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 16028 16532 16080 16584
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 11980 16396 12032 16448
rect 13268 16464 13320 16516
rect 12624 16439 12676 16448
rect 12624 16405 12641 16439
rect 12641 16405 12675 16439
rect 12675 16405 12676 16439
rect 12624 16396 12676 16405
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 13544 16396 13596 16448
rect 14556 16439 14608 16448
rect 14556 16405 14589 16439
rect 14589 16405 14608 16439
rect 14556 16396 14608 16405
rect 16856 16439 16908 16448
rect 16856 16405 16865 16439
rect 16865 16405 16899 16439
rect 16899 16405 16908 16439
rect 16856 16396 16908 16405
rect 3829 16294 3881 16346
rect 3893 16294 3945 16346
rect 3957 16294 4009 16346
rect 4021 16294 4073 16346
rect 4085 16294 4137 16346
rect 8268 16294 8320 16346
rect 8332 16294 8384 16346
rect 8396 16294 8448 16346
rect 8460 16294 8512 16346
rect 8524 16294 8576 16346
rect 12707 16294 12759 16346
rect 12771 16294 12823 16346
rect 12835 16294 12887 16346
rect 12899 16294 12951 16346
rect 12963 16294 13015 16346
rect 17146 16294 17198 16346
rect 17210 16294 17262 16346
rect 17274 16294 17326 16346
rect 17338 16294 17390 16346
rect 17402 16294 17454 16346
rect 5632 16192 5684 16244
rect 10600 16192 10652 16244
rect 4436 16124 4488 16176
rect 848 15988 900 16040
rect 2780 16099 2832 16108
rect 2780 16065 2789 16099
rect 2789 16065 2823 16099
rect 2823 16065 2832 16099
rect 2780 16056 2832 16065
rect 2964 16099 3016 16108
rect 2964 16065 2973 16099
rect 2973 16065 3007 16099
rect 3007 16065 3016 16099
rect 2964 16056 3016 16065
rect 2596 15988 2648 16040
rect 3240 15988 3292 16040
rect 9220 16124 9272 16176
rect 11796 16124 11848 16176
rect 12532 16192 12584 16244
rect 15384 16235 15436 16244
rect 15384 16201 15393 16235
rect 15393 16201 15427 16235
rect 15427 16201 15436 16235
rect 15384 16192 15436 16201
rect 15568 16235 15620 16244
rect 15568 16201 15577 16235
rect 15577 16201 15611 16235
rect 15611 16201 15620 16235
rect 15568 16192 15620 16201
rect 4712 16056 4764 16108
rect 5908 16056 5960 16108
rect 6460 16056 6512 16108
rect 8668 16099 8720 16108
rect 8668 16065 8672 16099
rect 8672 16065 8706 16099
rect 8706 16065 8720 16099
rect 8668 16056 8720 16065
rect 8760 16099 8812 16108
rect 8760 16065 8769 16099
rect 8769 16065 8803 16099
rect 8803 16065 8812 16099
rect 8760 16056 8812 16065
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 9036 16099 9088 16108
rect 6828 15988 6880 16040
rect 9036 16065 9044 16099
rect 9044 16065 9078 16099
rect 9078 16065 9088 16099
rect 9036 16056 9088 16065
rect 9128 16099 9180 16108
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 6920 15920 6972 15972
rect 5172 15852 5224 15904
rect 5448 15895 5500 15904
rect 5448 15861 5457 15895
rect 5457 15861 5491 15895
rect 5491 15861 5500 15895
rect 5448 15852 5500 15861
rect 5816 15895 5868 15904
rect 5816 15861 5825 15895
rect 5825 15861 5859 15895
rect 5859 15861 5868 15895
rect 5816 15852 5868 15861
rect 7380 15852 7432 15904
rect 7932 15852 7984 15904
rect 8208 15895 8260 15904
rect 8208 15861 8217 15895
rect 8217 15861 8251 15895
rect 8251 15861 8260 15895
rect 8208 15852 8260 15861
rect 8484 15963 8536 15972
rect 8484 15929 8493 15963
rect 8493 15929 8527 15963
rect 8527 15929 8536 15963
rect 8484 15920 8536 15929
rect 8760 15920 8812 15972
rect 11612 15988 11664 16040
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 13544 16056 13596 16108
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 12992 15988 13044 16040
rect 15476 16124 15528 16176
rect 16672 16192 16724 16244
rect 12532 15963 12584 15972
rect 12532 15929 12541 15963
rect 12541 15929 12575 15963
rect 12575 15929 12584 15963
rect 12532 15920 12584 15929
rect 17684 15988 17736 16040
rect 10324 15852 10376 15904
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 11704 15852 11756 15904
rect 11888 15852 11940 15904
rect 13084 15852 13136 15904
rect 3169 15750 3221 15802
rect 3233 15750 3285 15802
rect 3297 15750 3349 15802
rect 3361 15750 3413 15802
rect 3425 15750 3477 15802
rect 7608 15750 7660 15802
rect 7672 15750 7724 15802
rect 7736 15750 7788 15802
rect 7800 15750 7852 15802
rect 7864 15750 7916 15802
rect 12047 15750 12099 15802
rect 12111 15750 12163 15802
rect 12175 15750 12227 15802
rect 12239 15750 12291 15802
rect 12303 15750 12355 15802
rect 16486 15750 16538 15802
rect 16550 15750 16602 15802
rect 16614 15750 16666 15802
rect 16678 15750 16730 15802
rect 16742 15750 16794 15802
rect 2872 15648 2924 15700
rect 3516 15648 3568 15700
rect 5080 15691 5132 15700
rect 5080 15657 5089 15691
rect 5089 15657 5123 15691
rect 5123 15657 5132 15691
rect 5080 15648 5132 15657
rect 6920 15648 6972 15700
rect 10232 15580 10284 15632
rect 12992 15648 13044 15700
rect 1676 15512 1728 15564
rect 2596 15512 2648 15564
rect 6828 15555 6880 15564
rect 6828 15521 6837 15555
rect 6837 15521 6871 15555
rect 6871 15521 6880 15555
rect 6828 15512 6880 15521
rect 7288 15512 7340 15564
rect 7380 15512 7432 15564
rect 8300 15512 8352 15564
rect 11244 15512 11296 15564
rect 11888 15512 11940 15564
rect 11980 15512 12032 15564
rect 16856 15512 16908 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 1492 15444 1544 15496
rect 3608 15444 3660 15496
rect 5816 15444 5868 15496
rect 11336 15444 11388 15496
rect 12072 15487 12124 15496
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 2320 15376 2372 15428
rect 3332 15376 3384 15428
rect 940 15308 992 15360
rect 2412 15308 2464 15360
rect 3148 15308 3200 15360
rect 4252 15376 4304 15428
rect 11244 15376 11296 15428
rect 13084 15376 13136 15428
rect 16396 15376 16448 15428
rect 17776 15487 17828 15496
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 19248 15376 19300 15428
rect 4804 15308 4856 15360
rect 8300 15308 8352 15360
rect 8668 15308 8720 15360
rect 9956 15308 10008 15360
rect 10876 15308 10928 15360
rect 11612 15308 11664 15360
rect 14096 15308 14148 15360
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 15016 15351 15068 15360
rect 15016 15317 15025 15351
rect 15025 15317 15059 15351
rect 15059 15317 15068 15351
rect 15016 15308 15068 15317
rect 18328 15351 18380 15360
rect 18328 15317 18337 15351
rect 18337 15317 18371 15351
rect 18371 15317 18380 15351
rect 18328 15308 18380 15317
rect 3829 15206 3881 15258
rect 3893 15206 3945 15258
rect 3957 15206 4009 15258
rect 4021 15206 4073 15258
rect 4085 15206 4137 15258
rect 8268 15206 8320 15258
rect 8332 15206 8384 15258
rect 8396 15206 8448 15258
rect 8460 15206 8512 15258
rect 8524 15206 8576 15258
rect 12707 15206 12759 15258
rect 12771 15206 12823 15258
rect 12835 15206 12887 15258
rect 12899 15206 12951 15258
rect 12963 15206 13015 15258
rect 17146 15206 17198 15258
rect 17210 15206 17262 15258
rect 17274 15206 17326 15258
rect 17338 15206 17390 15258
rect 17402 15206 17454 15258
rect 2320 15104 2372 15156
rect 1492 14968 1544 15020
rect 2964 15104 3016 15156
rect 2780 15036 2832 15088
rect 6460 15104 6512 15156
rect 6828 15104 6880 15156
rect 4436 15036 4488 15088
rect 5724 15036 5776 15088
rect 6552 15036 6604 15088
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 2688 14943 2740 14952
rect 2688 14909 2697 14943
rect 2697 14909 2731 14943
rect 2731 14909 2740 14943
rect 2688 14900 2740 14909
rect 3332 14900 3384 14952
rect 4528 14968 4580 15020
rect 4988 15011 5040 15020
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 4436 14900 4488 14952
rect 2044 14832 2096 14884
rect 2412 14832 2464 14884
rect 5080 14832 5132 14884
rect 4068 14764 4120 14816
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 5356 14968 5408 15020
rect 6276 14968 6328 15020
rect 7288 15036 7340 15088
rect 8024 15147 8076 15156
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 8116 15104 8168 15156
rect 8392 15104 8444 15156
rect 9220 15104 9272 15156
rect 15292 15104 15344 15156
rect 16212 15104 16264 15156
rect 17776 15104 17828 15156
rect 5908 14900 5960 14952
rect 6920 14968 6972 15020
rect 10416 15036 10468 15088
rect 11428 15036 11480 15088
rect 12992 15036 13044 15088
rect 14280 15079 14332 15088
rect 14280 15045 14289 15079
rect 14289 15045 14323 15079
rect 14323 15045 14332 15079
rect 14280 15036 14332 15045
rect 16028 15036 16080 15088
rect 6460 14900 6512 14952
rect 6736 14832 6788 14884
rect 4620 14764 4672 14773
rect 5908 14807 5960 14816
rect 5908 14773 5917 14807
rect 5917 14773 5951 14807
rect 5951 14773 5960 14807
rect 5908 14764 5960 14773
rect 6460 14764 6512 14816
rect 7288 14900 7340 14952
rect 7472 14943 7524 14952
rect 7472 14909 7481 14943
rect 7481 14909 7515 14943
rect 7515 14909 7524 14943
rect 7472 14900 7524 14909
rect 8024 15011 8076 15020
rect 8024 14977 8033 15011
rect 8033 14977 8067 15011
rect 8067 14977 8076 15011
rect 8024 14968 8076 14977
rect 8300 14968 8352 15020
rect 8576 14968 8628 15020
rect 8852 15014 8904 15020
rect 8852 14980 8860 15014
rect 8860 14980 8894 15014
rect 8894 14980 8904 15014
rect 8852 14968 8904 14980
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 15292 14968 15344 15020
rect 8116 14900 8168 14952
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 10048 14900 10100 14952
rect 11888 14900 11940 14952
rect 10692 14832 10744 14884
rect 8484 14764 8536 14816
rect 9220 14764 9272 14816
rect 10508 14764 10560 14816
rect 16120 14900 16172 14952
rect 15016 14832 15068 14884
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 14648 14764 14700 14816
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 15936 14764 15988 14816
rect 3169 14662 3221 14714
rect 3233 14662 3285 14714
rect 3297 14662 3349 14714
rect 3361 14662 3413 14714
rect 3425 14662 3477 14714
rect 7608 14662 7660 14714
rect 7672 14662 7724 14714
rect 7736 14662 7788 14714
rect 7800 14662 7852 14714
rect 7864 14662 7916 14714
rect 12047 14662 12099 14714
rect 12111 14662 12163 14714
rect 12175 14662 12227 14714
rect 12239 14662 12291 14714
rect 12303 14662 12355 14714
rect 16486 14662 16538 14714
rect 16550 14662 16602 14714
rect 16614 14662 16666 14714
rect 16678 14662 16730 14714
rect 16742 14662 16794 14714
rect 1400 14560 1452 14612
rect 1952 14492 2004 14544
rect 4620 14560 4672 14612
rect 6184 14560 6236 14612
rect 7104 14560 7156 14612
rect 10968 14560 11020 14612
rect 11244 14560 11296 14612
rect 7380 14492 7432 14544
rect 1492 14424 1544 14476
rect 2964 14424 3016 14476
rect 1216 14356 1268 14408
rect 5724 14356 5776 14408
rect 6460 14399 6512 14408
rect 6460 14365 6469 14399
rect 6469 14365 6503 14399
rect 6503 14365 6512 14399
rect 6460 14356 6512 14365
rect 7564 14356 7616 14408
rect 8116 14356 8168 14408
rect 8760 14492 8812 14544
rect 8944 14492 8996 14544
rect 756 14288 808 14340
rect 3976 14288 4028 14340
rect 4160 14288 4212 14340
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 1676 14220 1728 14272
rect 4344 14220 4396 14272
rect 6828 14288 6880 14340
rect 9312 14467 9364 14476
rect 9312 14433 9321 14467
rect 9321 14433 9355 14467
rect 9355 14433 9364 14467
rect 9312 14424 9364 14433
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 10140 14424 10192 14476
rect 11888 14424 11940 14476
rect 13912 14492 13964 14544
rect 14372 14560 14424 14612
rect 15384 14492 15436 14544
rect 19064 14492 19116 14544
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 6920 14220 6972 14272
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 9588 14288 9640 14340
rect 9404 14220 9456 14272
rect 10140 14220 10192 14272
rect 13820 14356 13872 14408
rect 14372 14399 14424 14408
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 15568 14399 15620 14408
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 19156 14356 19208 14408
rect 12532 14220 12584 14272
rect 13360 14220 13412 14272
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 14280 14288 14332 14340
rect 16304 14288 16356 14340
rect 15660 14220 15712 14272
rect 15844 14220 15896 14272
rect 3829 14118 3881 14170
rect 3893 14118 3945 14170
rect 3957 14118 4009 14170
rect 4021 14118 4073 14170
rect 4085 14118 4137 14170
rect 8268 14118 8320 14170
rect 8332 14118 8384 14170
rect 8396 14118 8448 14170
rect 8460 14118 8512 14170
rect 8524 14118 8576 14170
rect 12707 14118 12759 14170
rect 12771 14118 12823 14170
rect 12835 14118 12887 14170
rect 12899 14118 12951 14170
rect 12963 14118 13015 14170
rect 17146 14118 17198 14170
rect 17210 14118 17262 14170
rect 17274 14118 17326 14170
rect 17338 14118 17390 14170
rect 17402 14118 17454 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 3056 13880 3108 13932
rect 3700 13948 3752 14000
rect 5356 14016 5408 14068
rect 8024 14016 8076 14068
rect 11336 14016 11388 14068
rect 12624 14016 12676 14068
rect 12992 14016 13044 14068
rect 13544 14016 13596 14068
rect 4160 13923 4212 13932
rect 4160 13889 4170 13923
rect 4170 13889 4204 13923
rect 4204 13889 4212 13923
rect 4160 13880 4212 13889
rect 4344 13923 4396 13932
rect 4344 13889 4353 13923
rect 4353 13889 4387 13923
rect 4387 13889 4396 13923
rect 4344 13880 4396 13889
rect 6092 13991 6144 14000
rect 6092 13957 6101 13991
rect 6101 13957 6135 13991
rect 6135 13957 6144 13991
rect 6092 13948 6144 13957
rect 6920 13948 6972 14000
rect 7104 13948 7156 14000
rect 9312 13948 9364 14000
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2872 13812 2924 13864
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 1952 13676 2004 13728
rect 2596 13676 2648 13728
rect 4896 13812 4948 13864
rect 7472 13880 7524 13932
rect 9404 13880 9456 13932
rect 9956 13948 10008 14000
rect 14004 14016 14056 14068
rect 16212 14016 16264 14068
rect 14096 13991 14148 14000
rect 14096 13957 14105 13991
rect 14105 13957 14139 13991
rect 14139 13957 14148 13991
rect 14096 13948 14148 13957
rect 14556 13948 14608 14000
rect 7012 13812 7064 13864
rect 8668 13812 8720 13864
rect 6092 13744 6144 13796
rect 7104 13744 7156 13796
rect 9220 13787 9272 13796
rect 9220 13753 9229 13787
rect 9229 13753 9263 13787
rect 9263 13753 9272 13787
rect 10232 13880 10284 13932
rect 10416 13880 10468 13932
rect 9680 13855 9732 13864
rect 9680 13821 9689 13855
rect 9689 13821 9723 13855
rect 9723 13821 9732 13855
rect 9680 13812 9732 13821
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 12532 13880 12584 13932
rect 12992 13880 13044 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 9772 13812 9824 13821
rect 13636 13812 13688 13864
rect 13912 13812 13964 13864
rect 14464 13812 14516 13864
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 15016 13812 15068 13864
rect 16304 13812 16356 13864
rect 9220 13744 9272 13753
rect 5172 13676 5224 13728
rect 7472 13676 7524 13728
rect 9312 13676 9364 13728
rect 10784 13744 10836 13796
rect 14280 13744 14332 13796
rect 11888 13676 11940 13728
rect 13084 13676 13136 13728
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 13728 13676 13780 13685
rect 3169 13574 3221 13626
rect 3233 13574 3285 13626
rect 3297 13574 3349 13626
rect 3361 13574 3413 13626
rect 3425 13574 3477 13626
rect 7608 13574 7660 13626
rect 7672 13574 7724 13626
rect 7736 13574 7788 13626
rect 7800 13574 7852 13626
rect 7864 13574 7916 13626
rect 12047 13574 12099 13626
rect 12111 13574 12163 13626
rect 12175 13574 12227 13626
rect 12239 13574 12291 13626
rect 12303 13574 12355 13626
rect 16486 13574 16538 13626
rect 16550 13574 16602 13626
rect 16614 13574 16666 13626
rect 16678 13574 16730 13626
rect 16742 13574 16794 13626
rect 2504 13472 2556 13524
rect 4068 13472 4120 13524
rect 4436 13472 4488 13524
rect 9956 13472 10008 13524
rect 10416 13472 10468 13524
rect 13268 13472 13320 13524
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 13728 13472 13780 13524
rect 13912 13472 13964 13524
rect 4160 13336 4212 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 1676 13268 1728 13320
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 1952 13311 2004 13320
rect 1952 13277 1961 13311
rect 1961 13277 1995 13311
rect 1995 13277 2004 13311
rect 1952 13268 2004 13277
rect 3148 13268 3200 13320
rect 3700 13268 3752 13320
rect 7472 13404 7524 13456
rect 8116 13404 8168 13456
rect 4528 13379 4580 13388
rect 4528 13345 4537 13379
rect 4537 13345 4571 13379
rect 4571 13345 4580 13379
rect 4528 13336 4580 13345
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 7656 13336 7708 13388
rect 8024 13336 8076 13388
rect 11888 13404 11940 13456
rect 12256 13404 12308 13456
rect 12900 13404 12952 13456
rect 15200 13472 15252 13524
rect 15384 13472 15436 13524
rect 16028 13472 16080 13524
rect 6736 13268 6788 13320
rect 9680 13268 9732 13320
rect 10876 13268 10928 13320
rect 10968 13268 11020 13320
rect 1768 13132 1820 13184
rect 1860 13132 1912 13184
rect 2320 13132 2372 13184
rect 2412 13132 2464 13184
rect 2596 13132 2648 13184
rect 3608 13243 3660 13252
rect 3608 13209 3617 13243
rect 3617 13209 3651 13243
rect 3651 13209 3660 13243
rect 3608 13200 3660 13209
rect 4712 13200 4764 13252
rect 5724 13200 5776 13252
rect 6000 13243 6052 13252
rect 6000 13209 6009 13243
rect 6009 13209 6043 13243
rect 6043 13209 6052 13243
rect 6000 13200 6052 13209
rect 6092 13200 6144 13252
rect 10140 13200 10192 13252
rect 11244 13243 11296 13252
rect 11244 13209 11253 13243
rect 11253 13209 11287 13243
rect 11287 13209 11296 13243
rect 11244 13200 11296 13209
rect 11336 13200 11388 13252
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12256 13311 12308 13320
rect 12256 13277 12265 13311
rect 12265 13277 12299 13311
rect 12299 13277 12308 13311
rect 12256 13268 12308 13277
rect 14740 13379 14792 13388
rect 14740 13345 14749 13379
rect 14749 13345 14783 13379
rect 14783 13345 14792 13379
rect 14740 13336 14792 13345
rect 15016 13336 15068 13388
rect 15384 13379 15436 13388
rect 15384 13345 15393 13379
rect 15393 13345 15427 13379
rect 15427 13345 15436 13379
rect 15384 13336 15436 13345
rect 13452 13268 13504 13320
rect 15292 13311 15344 13320
rect 15292 13277 15300 13311
rect 15300 13277 15334 13311
rect 15334 13277 15344 13311
rect 15292 13268 15344 13277
rect 18604 13404 18656 13456
rect 15752 13336 15804 13388
rect 13544 13200 13596 13252
rect 14096 13200 14148 13252
rect 14280 13200 14332 13252
rect 5080 13132 5132 13184
rect 5632 13132 5684 13184
rect 6736 13132 6788 13184
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 9404 13132 9456 13184
rect 9772 13132 9824 13184
rect 11888 13132 11940 13184
rect 13452 13132 13504 13184
rect 14924 13132 14976 13184
rect 16488 13268 16540 13320
rect 16672 13243 16724 13252
rect 16672 13209 16681 13243
rect 16681 13209 16715 13243
rect 16715 13209 16724 13243
rect 16672 13200 16724 13209
rect 17592 13132 17644 13184
rect 3829 13030 3881 13082
rect 3893 13030 3945 13082
rect 3957 13030 4009 13082
rect 4021 13030 4073 13082
rect 4085 13030 4137 13082
rect 8268 13030 8320 13082
rect 8332 13030 8384 13082
rect 8396 13030 8448 13082
rect 8460 13030 8512 13082
rect 8524 13030 8576 13082
rect 12707 13030 12759 13082
rect 12771 13030 12823 13082
rect 12835 13030 12887 13082
rect 12899 13030 12951 13082
rect 12963 13030 13015 13082
rect 17146 13030 17198 13082
rect 17210 13030 17262 13082
rect 17274 13030 17326 13082
rect 17338 13030 17390 13082
rect 17402 13030 17454 13082
rect 2964 12928 3016 12980
rect 3424 12928 3476 12980
rect 3792 12928 3844 12980
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 2688 12792 2740 12844
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 1032 12588 1084 12640
rect 7656 12860 7708 12912
rect 9128 12928 9180 12980
rect 5172 12792 5224 12844
rect 3700 12588 3752 12640
rect 4160 12588 4212 12640
rect 4620 12588 4672 12640
rect 6184 12792 6236 12844
rect 6460 12792 6512 12844
rect 8300 12835 8352 12844
rect 8300 12801 8304 12835
rect 8304 12801 8338 12835
rect 8338 12801 8352 12835
rect 8300 12792 8352 12801
rect 8852 12860 8904 12912
rect 8944 12860 8996 12912
rect 10416 12928 10468 12980
rect 11152 12928 11204 12980
rect 12164 12928 12216 12980
rect 12256 12928 12308 12980
rect 12808 12928 12860 12980
rect 7472 12724 7524 12776
rect 9680 12792 9732 12844
rect 10876 12860 10928 12912
rect 13728 12928 13780 12980
rect 14188 12928 14240 12980
rect 13636 12860 13688 12912
rect 15476 12928 15528 12980
rect 15844 12928 15896 12980
rect 16396 12928 16448 12980
rect 15200 12860 15252 12912
rect 17040 12928 17092 12980
rect 19340 12860 19392 12912
rect 9496 12724 9548 12776
rect 9864 12767 9916 12776
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 9864 12724 9916 12733
rect 5724 12588 5776 12640
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 7932 12588 7984 12640
rect 8024 12588 8076 12640
rect 8852 12656 8904 12708
rect 11704 12724 11756 12776
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 14004 12835 14056 12844
rect 14004 12801 14013 12835
rect 14013 12801 14047 12835
rect 14047 12801 14056 12835
rect 14004 12792 14056 12801
rect 10048 12656 10100 12708
rect 11152 12656 11204 12708
rect 13912 12724 13964 12776
rect 14832 12792 14884 12844
rect 15108 12792 15160 12844
rect 15016 12724 15068 12776
rect 15844 12792 15896 12844
rect 16028 12835 16080 12844
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 16672 12792 16724 12844
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 17500 12835 17552 12844
rect 17500 12801 17509 12835
rect 17509 12801 17543 12835
rect 17543 12801 17552 12835
rect 17500 12792 17552 12801
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 16396 12724 16448 12776
rect 15568 12699 15620 12708
rect 15568 12665 15577 12699
rect 15577 12665 15611 12699
rect 15611 12665 15620 12699
rect 15568 12656 15620 12665
rect 9864 12588 9916 12640
rect 13544 12588 13596 12640
rect 13820 12588 13872 12640
rect 15292 12588 15344 12640
rect 15752 12588 15804 12640
rect 3169 12486 3221 12538
rect 3233 12486 3285 12538
rect 3297 12486 3349 12538
rect 3361 12486 3413 12538
rect 3425 12486 3477 12538
rect 7608 12486 7660 12538
rect 7672 12486 7724 12538
rect 7736 12486 7788 12538
rect 7800 12486 7852 12538
rect 7864 12486 7916 12538
rect 12047 12486 12099 12538
rect 12111 12486 12163 12538
rect 12175 12486 12227 12538
rect 12239 12486 12291 12538
rect 12303 12486 12355 12538
rect 16486 12486 16538 12538
rect 16550 12486 16602 12538
rect 16614 12486 16666 12538
rect 16678 12486 16730 12538
rect 16742 12486 16794 12538
rect 3608 12384 3660 12436
rect 4160 12384 4212 12436
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 1860 12316 1912 12368
rect 7748 12384 7800 12436
rect 8300 12384 8352 12436
rect 9404 12384 9456 12436
rect 9864 12384 9916 12436
rect 11244 12384 11296 12436
rect 11796 12384 11848 12436
rect 13912 12384 13964 12436
rect 14464 12384 14516 12436
rect 15660 12384 15712 12436
rect 6644 12316 6696 12368
rect 7288 12316 7340 12368
rect 848 12248 900 12300
rect 1216 12248 1268 12300
rect 1124 12180 1176 12232
rect 1584 12155 1636 12164
rect 1584 12121 1593 12155
rect 1593 12121 1627 12155
rect 1627 12121 1636 12155
rect 1584 12112 1636 12121
rect 2044 12180 2096 12232
rect 2596 12248 2648 12300
rect 4252 12223 4304 12232
rect 4252 12189 4261 12223
rect 4261 12189 4295 12223
rect 4295 12189 4304 12223
rect 4252 12180 4304 12189
rect 3148 12112 3200 12164
rect 5540 12248 5592 12300
rect 6000 12248 6052 12300
rect 7748 12248 7800 12300
rect 5356 12180 5408 12232
rect 7012 12180 7064 12232
rect 14096 12316 14148 12368
rect 11704 12248 11756 12300
rect 12624 12248 12676 12300
rect 13912 12248 13964 12300
rect 15936 12291 15988 12300
rect 15936 12257 15945 12291
rect 15945 12257 15979 12291
rect 15979 12257 15988 12291
rect 15936 12248 15988 12257
rect 9128 12180 9180 12232
rect 9496 12180 9548 12232
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 14832 12180 14884 12232
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 5816 12112 5868 12164
rect 7196 12112 7248 12164
rect 7472 12112 7524 12164
rect 7748 12155 7800 12164
rect 7748 12121 7757 12155
rect 7757 12121 7791 12155
rect 7791 12121 7800 12155
rect 7748 12112 7800 12121
rect 8116 12112 8168 12164
rect 8484 12112 8536 12164
rect 13268 12112 13320 12164
rect 1676 12044 1728 12096
rect 2872 12044 2924 12096
rect 4344 12044 4396 12096
rect 5172 12044 5224 12096
rect 6276 12044 6328 12096
rect 6552 12044 6604 12096
rect 8760 12044 8812 12096
rect 9588 12044 9640 12096
rect 10416 12044 10468 12096
rect 11060 12044 11112 12096
rect 11704 12044 11756 12096
rect 15476 12112 15528 12164
rect 14188 12044 14240 12096
rect 14464 12044 14516 12096
rect 15292 12044 15344 12096
rect 3829 11942 3881 11994
rect 3893 11942 3945 11994
rect 3957 11942 4009 11994
rect 4021 11942 4073 11994
rect 4085 11942 4137 11994
rect 8268 11942 8320 11994
rect 8332 11942 8384 11994
rect 8396 11942 8448 11994
rect 8460 11942 8512 11994
rect 8524 11942 8576 11994
rect 12707 11942 12759 11994
rect 12771 11942 12823 11994
rect 12835 11942 12887 11994
rect 12899 11942 12951 11994
rect 12963 11942 13015 11994
rect 17146 11942 17198 11994
rect 17210 11942 17262 11994
rect 17274 11942 17326 11994
rect 17338 11942 17390 11994
rect 17402 11942 17454 11994
rect 572 11840 624 11892
rect 2872 11772 2924 11824
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 2136 11704 2188 11756
rect 2412 11747 2464 11756
rect 2412 11713 2416 11747
rect 2416 11713 2450 11747
rect 2450 11713 2464 11747
rect 2412 11704 2464 11713
rect 1952 11636 2004 11688
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 3700 11772 3752 11824
rect 4068 11772 4120 11824
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 4620 11704 4672 11756
rect 5356 11704 5408 11756
rect 7104 11840 7156 11892
rect 7932 11883 7984 11892
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 8024 11840 8076 11892
rect 9220 11840 9272 11892
rect 9404 11840 9456 11892
rect 13912 11840 13964 11892
rect 15476 11840 15528 11892
rect 16396 11840 16448 11892
rect 16856 11840 16908 11892
rect 2504 11568 2556 11620
rect 2780 11568 2832 11620
rect 1584 11500 1636 11552
rect 1860 11500 1912 11552
rect 3148 11500 3200 11552
rect 5540 11636 5592 11688
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 8852 11772 8904 11824
rect 11336 11772 11388 11824
rect 16304 11772 16356 11824
rect 16488 11772 16540 11824
rect 9220 11704 9272 11756
rect 10968 11704 11020 11756
rect 11796 11704 11848 11756
rect 4712 11568 4764 11620
rect 5264 11568 5316 11620
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 7656 11636 7708 11688
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 8576 11636 8628 11688
rect 13084 11636 13136 11688
rect 13728 11704 13780 11756
rect 14188 11704 14240 11756
rect 14740 11704 14792 11756
rect 17316 11772 17368 11824
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 5356 11500 5408 11552
rect 6092 11500 6144 11552
rect 6828 11500 6880 11552
rect 11060 11568 11112 11620
rect 8576 11500 8628 11552
rect 9220 11500 9272 11552
rect 9312 11500 9364 11552
rect 12900 11568 12952 11620
rect 14464 11636 14516 11688
rect 11336 11500 11388 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 16028 11500 16080 11552
rect 18144 11636 18196 11688
rect 17500 11568 17552 11620
rect 18420 11500 18472 11552
rect 3169 11398 3221 11450
rect 3233 11398 3285 11450
rect 3297 11398 3349 11450
rect 3361 11398 3413 11450
rect 3425 11398 3477 11450
rect 7608 11398 7660 11450
rect 7672 11398 7724 11450
rect 7736 11398 7788 11450
rect 7800 11398 7852 11450
rect 7864 11398 7916 11450
rect 12047 11398 12099 11450
rect 12111 11398 12163 11450
rect 12175 11398 12227 11450
rect 12239 11398 12291 11450
rect 12303 11398 12355 11450
rect 16486 11398 16538 11450
rect 16550 11398 16602 11450
rect 16614 11398 16666 11450
rect 16678 11398 16730 11450
rect 16742 11398 16794 11450
rect 4620 11296 4672 11348
rect 5816 11339 5868 11348
rect 5816 11305 5825 11339
rect 5825 11305 5859 11339
rect 5859 11305 5868 11339
rect 5816 11296 5868 11305
rect 6828 11296 6880 11348
rect 7288 11296 7340 11348
rect 7564 11296 7616 11348
rect 1308 11228 1360 11280
rect 3976 11228 4028 11280
rect 6000 11228 6052 11280
rect 6276 11228 6328 11280
rect 11336 11296 11388 11348
rect 11520 11296 11572 11348
rect 15016 11296 15068 11348
rect 15292 11296 15344 11348
rect 15936 11339 15988 11348
rect 15936 11305 15945 11339
rect 15945 11305 15979 11339
rect 15979 11305 15988 11339
rect 15936 11296 15988 11305
rect 2596 11160 2648 11212
rect 4160 11160 4212 11212
rect 6552 11160 6604 11212
rect 9036 11228 9088 11280
rect 9404 11228 9456 11280
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2044 11092 2096 11144
rect 4528 11092 4580 11144
rect 6000 11092 6052 11144
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 9496 11160 9548 11212
rect 13728 11160 13780 11212
rect 1676 11024 1728 11076
rect 1952 11024 2004 11076
rect 2688 11024 2740 11076
rect 5264 11024 5316 11076
rect 5724 11024 5776 11076
rect 7288 11067 7340 11076
rect 7288 11033 7297 11067
rect 7297 11033 7331 11067
rect 7331 11033 7340 11067
rect 7288 11024 7340 11033
rect 7564 11024 7616 11076
rect 9312 11092 9364 11144
rect 9772 11092 9824 11144
rect 12164 11092 12216 11144
rect 12624 11092 12676 11144
rect 13636 11092 13688 11144
rect 16028 11228 16080 11280
rect 16672 11228 16724 11280
rect 17868 11228 17920 11280
rect 9588 11024 9640 11076
rect 13452 11024 13504 11076
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 3424 10956 3476 11008
rect 4068 10956 4120 11008
rect 6552 10956 6604 11008
rect 7932 10956 7984 11008
rect 8116 10956 8168 11008
rect 11060 10956 11112 11008
rect 13728 11067 13780 11076
rect 13728 11033 13737 11067
rect 13737 11033 13771 11067
rect 13771 11033 13780 11067
rect 13728 11024 13780 11033
rect 14556 11135 14608 11144
rect 14556 11101 14565 11135
rect 14565 11101 14599 11135
rect 14599 11101 14608 11135
rect 14556 11092 14608 11101
rect 14648 11092 14700 11144
rect 14924 11135 14976 11144
rect 14924 11101 14933 11135
rect 14933 11101 14967 11135
rect 14967 11101 14976 11135
rect 14924 11092 14976 11101
rect 16396 11092 16448 11144
rect 15752 11024 15804 11076
rect 16580 11135 16632 11144
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 16948 11092 17000 11144
rect 18420 11092 18472 11144
rect 17316 11067 17368 11076
rect 17316 11033 17325 11067
rect 17325 11033 17359 11067
rect 17359 11033 17368 11067
rect 17316 11024 17368 11033
rect 17868 11024 17920 11076
rect 13912 10956 13964 11008
rect 14832 10956 14884 11008
rect 15200 10956 15252 11008
rect 16120 10956 16172 11008
rect 3829 10854 3881 10906
rect 3893 10854 3945 10906
rect 3957 10854 4009 10906
rect 4021 10854 4073 10906
rect 4085 10854 4137 10906
rect 8268 10854 8320 10906
rect 8332 10854 8384 10906
rect 8396 10854 8448 10906
rect 8460 10854 8512 10906
rect 8524 10854 8576 10906
rect 12707 10854 12759 10906
rect 12771 10854 12823 10906
rect 12835 10854 12887 10906
rect 12899 10854 12951 10906
rect 12963 10854 13015 10906
rect 17146 10854 17198 10906
rect 17210 10854 17262 10906
rect 17274 10854 17326 10906
rect 17338 10854 17390 10906
rect 17402 10854 17454 10906
rect 2228 10752 2280 10804
rect 2412 10752 2464 10804
rect 3332 10752 3384 10804
rect 4620 10752 4672 10804
rect 4804 10752 4856 10804
rect 5264 10752 5316 10804
rect 5448 10752 5500 10804
rect 6460 10752 6512 10804
rect 6644 10752 6696 10804
rect 7472 10752 7524 10804
rect 7748 10752 7800 10804
rect 9404 10752 9456 10804
rect 1584 10684 1636 10736
rect 1952 10684 2004 10736
rect 5724 10684 5776 10736
rect 6368 10684 6420 10736
rect 7104 10727 7156 10736
rect 7104 10693 7113 10727
rect 7113 10693 7147 10727
rect 7147 10693 7156 10727
rect 7104 10684 7156 10693
rect 7380 10684 7432 10736
rect 7656 10684 7708 10736
rect 7840 10684 7892 10736
rect 8208 10684 8260 10736
rect 9588 10752 9640 10804
rect 10784 10752 10836 10804
rect 11244 10795 11296 10804
rect 11244 10761 11253 10795
rect 11253 10761 11287 10795
rect 11287 10761 11296 10795
rect 11244 10752 11296 10761
rect 12624 10752 12676 10804
rect 13544 10752 13596 10804
rect 16764 10752 16816 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 2872 10616 2924 10668
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 6736 10616 6788 10668
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 2136 10591 2188 10600
rect 2136 10557 2145 10591
rect 2145 10557 2179 10591
rect 2179 10557 2188 10591
rect 2136 10548 2188 10557
rect 3424 10591 3476 10600
rect 3424 10557 3433 10591
rect 3433 10557 3467 10591
rect 3467 10557 3476 10591
rect 3424 10548 3476 10557
rect 3976 10548 4028 10600
rect 5172 10548 5224 10600
rect 7104 10548 7156 10600
rect 11336 10684 11388 10736
rect 11888 10727 11940 10736
rect 11888 10693 11897 10727
rect 11897 10693 11931 10727
rect 11931 10693 11940 10727
rect 11888 10684 11940 10693
rect 9588 10616 9640 10668
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 14556 10684 14608 10736
rect 14648 10684 14700 10736
rect 17592 10684 17644 10736
rect 18880 10684 18932 10736
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 13544 10616 13596 10668
rect 16488 10616 16540 10668
rect 16672 10616 16724 10668
rect 17408 10616 17460 10668
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 18420 10616 18472 10668
rect 1584 10523 1636 10532
rect 1584 10489 1593 10523
rect 1593 10489 1627 10523
rect 1627 10489 1636 10523
rect 1584 10480 1636 10489
rect 4068 10523 4120 10532
rect 4068 10489 4077 10523
rect 4077 10489 4111 10523
rect 4111 10489 4120 10523
rect 4068 10480 4120 10489
rect 2320 10412 2372 10464
rect 2872 10412 2924 10464
rect 5908 10412 5960 10464
rect 7104 10412 7156 10464
rect 7656 10412 7708 10464
rect 8116 10412 8168 10464
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 8484 10523 8536 10532
rect 8484 10489 8493 10523
rect 8493 10489 8527 10523
rect 8527 10489 8536 10523
rect 8484 10480 8536 10489
rect 10232 10591 10284 10600
rect 10232 10557 10241 10591
rect 10241 10557 10275 10591
rect 10275 10557 10284 10591
rect 10232 10548 10284 10557
rect 11520 10548 11572 10600
rect 11980 10548 12032 10600
rect 12164 10548 12216 10600
rect 12992 10548 13044 10600
rect 13452 10548 13504 10600
rect 12624 10480 12676 10532
rect 14188 10480 14240 10532
rect 17040 10480 17092 10532
rect 10048 10412 10100 10464
rect 10232 10412 10284 10464
rect 11704 10412 11756 10464
rect 14648 10412 14700 10464
rect 14740 10412 14792 10464
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 16212 10412 16264 10464
rect 3169 10310 3221 10362
rect 3233 10310 3285 10362
rect 3297 10310 3349 10362
rect 3361 10310 3413 10362
rect 3425 10310 3477 10362
rect 7608 10310 7660 10362
rect 7672 10310 7724 10362
rect 7736 10310 7788 10362
rect 7800 10310 7852 10362
rect 7864 10310 7916 10362
rect 12047 10310 12099 10362
rect 12111 10310 12163 10362
rect 12175 10310 12227 10362
rect 12239 10310 12291 10362
rect 12303 10310 12355 10362
rect 16486 10310 16538 10362
rect 16550 10310 16602 10362
rect 16614 10310 16666 10362
rect 16678 10310 16730 10362
rect 16742 10310 16794 10362
rect 1400 10208 1452 10260
rect 1952 10140 2004 10192
rect 2136 10140 2188 10192
rect 4804 10208 4856 10260
rect 5448 10208 5500 10260
rect 5540 10208 5592 10260
rect 5908 10208 5960 10260
rect 3700 10140 3752 10192
rect 6644 10208 6696 10260
rect 7748 10208 7800 10260
rect 8208 10208 8260 10260
rect 8576 10208 8628 10260
rect 1860 10072 1912 10124
rect 2964 10072 3016 10124
rect 7196 10140 7248 10192
rect 8852 10140 8904 10192
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 9680 10208 9732 10260
rect 11980 10208 12032 10260
rect 9404 10140 9456 10192
rect 10784 10183 10836 10192
rect 10784 10149 10793 10183
rect 10793 10149 10827 10183
rect 10827 10149 10836 10183
rect 10784 10140 10836 10149
rect 11060 10140 11112 10192
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 15752 10208 15804 10260
rect 16028 10208 16080 10260
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 1952 10047 2004 10056
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 2136 10004 2188 10056
rect 4160 10004 4212 10056
rect 4528 10004 4580 10056
rect 2412 9936 2464 9988
rect 2688 9936 2740 9988
rect 3056 9936 3108 9988
rect 6276 10072 6328 10124
rect 6552 10072 6604 10124
rect 7288 10072 7340 10124
rect 5540 10004 5592 10056
rect 6184 10004 6236 10056
rect 7380 10004 7432 10056
rect 8208 10004 8260 10056
rect 9312 10004 9364 10056
rect 12164 10072 12216 10124
rect 4988 9936 5040 9988
rect 9680 9936 9732 9988
rect 10968 9936 11020 9988
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 11612 10004 11664 10056
rect 11980 10004 12032 10056
rect 14832 10072 14884 10124
rect 14924 10072 14976 10124
rect 13176 10004 13228 10056
rect 14648 10004 14700 10056
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 19432 10072 19484 10124
rect 3608 9868 3660 9920
rect 3792 9868 3844 9920
rect 3976 9868 4028 9920
rect 4712 9868 4764 9920
rect 5448 9868 5500 9920
rect 5540 9911 5592 9920
rect 5540 9877 5549 9911
rect 5549 9877 5583 9911
rect 5583 9877 5592 9911
rect 5540 9868 5592 9877
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 9588 9868 9640 9920
rect 10876 9868 10928 9920
rect 11244 9868 11296 9920
rect 13452 9936 13504 9988
rect 14464 9936 14516 9988
rect 16856 9936 16908 9988
rect 12348 9868 12400 9920
rect 13268 9868 13320 9920
rect 16212 9868 16264 9920
rect 17408 10004 17460 10056
rect 17960 10047 18012 10056
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 3829 9766 3881 9818
rect 3893 9766 3945 9818
rect 3957 9766 4009 9818
rect 4021 9766 4073 9818
rect 4085 9766 4137 9818
rect 8268 9766 8320 9818
rect 8332 9766 8384 9818
rect 8396 9766 8448 9818
rect 8460 9766 8512 9818
rect 8524 9766 8576 9818
rect 12707 9766 12759 9818
rect 12771 9766 12823 9818
rect 12835 9766 12887 9818
rect 12899 9766 12951 9818
rect 12963 9766 13015 9818
rect 17146 9766 17198 9818
rect 17210 9766 17262 9818
rect 17274 9766 17326 9818
rect 17338 9766 17390 9818
rect 17402 9766 17454 9818
rect 2044 9664 2096 9716
rect 1768 9596 1820 9648
rect 2688 9596 2740 9648
rect 3608 9664 3660 9716
rect 3792 9664 3844 9716
rect 7104 9664 7156 9716
rect 7472 9664 7524 9716
rect 5632 9596 5684 9648
rect 6552 9596 6604 9648
rect 7564 9596 7616 9648
rect 8208 9596 8260 9648
rect 9404 9664 9456 9716
rect 9680 9664 9732 9716
rect 10232 9664 10284 9716
rect 10692 9664 10744 9716
rect 10968 9664 11020 9716
rect 10508 9596 10560 9648
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 4068 9528 4120 9580
rect 4528 9460 4580 9512
rect 4988 9528 5040 9580
rect 6184 9528 6236 9580
rect 7104 9528 7156 9580
rect 9312 9528 9364 9580
rect 9680 9528 9732 9580
rect 13268 9664 13320 9716
rect 11244 9596 11296 9648
rect 6644 9460 6696 9512
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 8668 9460 8720 9512
rect 8852 9460 8904 9512
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 10508 9460 10560 9512
rect 4988 9392 5040 9444
rect 9680 9392 9732 9444
rect 11796 9596 11848 9648
rect 12992 9596 13044 9648
rect 11612 9528 11664 9580
rect 13636 9571 13688 9604
rect 13636 9552 13645 9571
rect 13645 9552 13679 9571
rect 13679 9552 13688 9571
rect 13268 9460 13320 9512
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 14096 9707 14148 9716
rect 14096 9673 14105 9707
rect 14105 9673 14139 9707
rect 14139 9673 14148 9707
rect 14096 9664 14148 9673
rect 14372 9664 14424 9716
rect 13912 9528 13964 9580
rect 14004 9528 14056 9580
rect 14096 9503 14148 9512
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 16028 9664 16080 9716
rect 16212 9664 16264 9716
rect 17960 9664 18012 9716
rect 16304 9596 16356 9648
rect 16948 9528 17000 9580
rect 15660 9460 15712 9512
rect 16304 9460 16356 9512
rect 16488 9460 16540 9512
rect 17316 9503 17368 9512
rect 17316 9469 17325 9503
rect 17325 9469 17359 9503
rect 17359 9469 17368 9503
rect 17316 9460 17368 9469
rect 3516 9324 3568 9376
rect 4528 9324 4580 9376
rect 6644 9324 6696 9376
rect 7104 9324 7156 9376
rect 8208 9324 8260 9376
rect 9588 9324 9640 9376
rect 15936 9392 15988 9444
rect 10508 9324 10560 9376
rect 11060 9324 11112 9376
rect 11796 9324 11848 9376
rect 11980 9324 12032 9376
rect 13084 9324 13136 9376
rect 14372 9324 14424 9376
rect 15384 9324 15436 9376
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16212 9324 16264 9333
rect 16764 9324 16816 9376
rect 17040 9324 17092 9376
rect 17132 9324 17184 9376
rect 18420 9528 18472 9580
rect 17868 9460 17920 9512
rect 18512 9324 18564 9376
rect 3169 9222 3221 9274
rect 3233 9222 3285 9274
rect 3297 9222 3349 9274
rect 3361 9222 3413 9274
rect 3425 9222 3477 9274
rect 7608 9222 7660 9274
rect 7672 9222 7724 9274
rect 7736 9222 7788 9274
rect 7800 9222 7852 9274
rect 7864 9222 7916 9274
rect 12047 9222 12099 9274
rect 12111 9222 12163 9274
rect 12175 9222 12227 9274
rect 12239 9222 12291 9274
rect 12303 9222 12355 9274
rect 16486 9222 16538 9274
rect 16550 9222 16602 9274
rect 16614 9222 16666 9274
rect 16678 9222 16730 9274
rect 16742 9222 16794 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 2596 9120 2648 9172
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3792 9120 3844 9172
rect 4160 9120 4212 9172
rect 4344 9120 4396 9172
rect 5448 9120 5500 9172
rect 6092 9120 6144 9172
rect 6920 9120 6972 9172
rect 7748 9120 7800 9172
rect 2228 9052 2280 9104
rect 3608 9052 3660 9104
rect 7012 9052 7064 9104
rect 9680 9120 9732 9172
rect 10324 9163 10376 9172
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 10692 9120 10744 9172
rect 13820 9120 13872 9172
rect 14832 9120 14884 9172
rect 15384 9120 15436 9172
rect 15660 9120 15712 9172
rect 16028 9120 16080 9172
rect 10968 9095 11020 9104
rect 10968 9061 10977 9095
rect 10977 9061 11011 9095
rect 11011 9061 11020 9095
rect 10968 9052 11020 9061
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2228 8916 2280 8968
rect 2872 8984 2924 9036
rect 5632 8984 5684 9036
rect 6920 8984 6972 9036
rect 7840 8984 7892 9036
rect 8392 8984 8444 9036
rect 10692 8984 10744 9036
rect 3240 8916 3292 8968
rect 4436 8916 4488 8968
rect 5448 8916 5500 8968
rect 2044 8848 2096 8900
rect 3056 8780 3108 8832
rect 4528 8780 4580 8832
rect 5632 8848 5684 8900
rect 7104 8916 7156 8968
rect 8760 8959 8812 8968
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9588 8959 9640 8968
rect 9588 8925 9597 8959
rect 9597 8925 9631 8959
rect 9631 8925 9640 8959
rect 9588 8916 9640 8925
rect 9772 8916 9824 8968
rect 10140 8916 10192 8968
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 11520 9052 11572 9104
rect 17316 9120 17368 9172
rect 7196 8848 7248 8900
rect 8208 8848 8260 8900
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 13544 8984 13596 9036
rect 16396 9052 16448 9104
rect 16764 8984 16816 9036
rect 17960 8984 18012 9036
rect 11612 8916 11664 8968
rect 12624 8916 12676 8968
rect 13636 8916 13688 8968
rect 13820 8916 13872 8968
rect 15016 8916 15068 8968
rect 16304 8916 16356 8968
rect 16396 8959 16448 8968
rect 16396 8925 16405 8959
rect 16405 8925 16439 8959
rect 16439 8925 16448 8959
rect 16396 8916 16448 8925
rect 11796 8848 11848 8900
rect 11612 8780 11664 8832
rect 12624 8780 12676 8832
rect 15108 8848 15160 8900
rect 15476 8848 15528 8900
rect 16028 8848 16080 8900
rect 14188 8780 14240 8832
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 14924 8780 14976 8832
rect 16304 8780 16356 8832
rect 17040 8848 17092 8900
rect 17408 8780 17460 8832
rect 3829 8678 3881 8730
rect 3893 8678 3945 8730
rect 3957 8678 4009 8730
rect 4021 8678 4073 8730
rect 4085 8678 4137 8730
rect 8268 8678 8320 8730
rect 8332 8678 8384 8730
rect 8396 8678 8448 8730
rect 8460 8678 8512 8730
rect 8524 8678 8576 8730
rect 12707 8678 12759 8730
rect 12771 8678 12823 8730
rect 12835 8678 12887 8730
rect 12899 8678 12951 8730
rect 12963 8678 13015 8730
rect 17146 8678 17198 8730
rect 17210 8678 17262 8730
rect 17274 8678 17326 8730
rect 17338 8678 17390 8730
rect 17402 8678 17454 8730
rect 2964 8576 3016 8628
rect 3516 8576 3568 8628
rect 3148 8508 3200 8560
rect 3608 8508 3660 8560
rect 5632 8508 5684 8560
rect 3700 8440 3752 8492
rect 6000 8576 6052 8628
rect 8392 8576 8444 8628
rect 9496 8576 9548 8628
rect 9588 8576 9640 8628
rect 10416 8576 10468 8628
rect 11612 8576 11664 8628
rect 12440 8576 12492 8628
rect 14004 8619 14056 8628
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 15844 8619 15896 8628
rect 15844 8585 15853 8619
rect 15853 8585 15887 8619
rect 15887 8585 15896 8619
rect 15844 8576 15896 8585
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 16948 8576 17000 8628
rect 17132 8576 17184 8628
rect 17224 8576 17276 8628
rect 17684 8576 17736 8628
rect 18420 8619 18472 8628
rect 18420 8585 18429 8619
rect 18429 8585 18463 8619
rect 18463 8585 18472 8619
rect 18420 8576 18472 8585
rect 7012 8508 7064 8560
rect 7564 8508 7616 8560
rect 8116 8551 8168 8560
rect 8116 8517 8125 8551
rect 8125 8517 8159 8551
rect 8159 8517 8168 8551
rect 8116 8508 8168 8517
rect 8484 8508 8536 8560
rect 8852 8508 8904 8560
rect 11152 8508 11204 8560
rect 11796 8508 11848 8560
rect 7196 8440 7248 8492
rect 8760 8440 8812 8492
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 10692 8440 10744 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 1216 8304 1268 8356
rect 8668 8372 8720 8424
rect 8852 8372 8904 8424
rect 15384 8508 15436 8560
rect 12900 8440 12952 8492
rect 12532 8372 12584 8424
rect 12624 8372 12676 8424
rect 13636 8372 13688 8424
rect 14188 8372 14240 8424
rect 16764 8440 16816 8492
rect 17224 8440 17276 8492
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 16396 8415 16448 8424
rect 6092 8304 6144 8356
rect 8484 8304 8536 8356
rect 8576 8304 8628 8356
rect 9036 8304 9088 8356
rect 11060 8304 11112 8356
rect 13544 8304 13596 8356
rect 15384 8347 15436 8356
rect 15384 8313 15393 8347
rect 15393 8313 15427 8347
rect 15427 8313 15436 8347
rect 15384 8304 15436 8313
rect 16396 8381 16405 8415
rect 16405 8381 16439 8415
rect 16439 8381 16448 8415
rect 16396 8372 16448 8381
rect 16948 8372 17000 8424
rect 17316 8415 17368 8424
rect 17316 8381 17325 8415
rect 17325 8381 17359 8415
rect 17359 8381 17368 8415
rect 17316 8372 17368 8381
rect 17684 8440 17736 8492
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 17960 8440 18012 8492
rect 17500 8415 17552 8424
rect 17500 8381 17509 8415
rect 17509 8381 17543 8415
rect 17543 8381 17552 8415
rect 17500 8372 17552 8381
rect 18512 8372 18564 8424
rect 1860 8236 1912 8288
rect 2964 8236 3016 8288
rect 3240 8236 3292 8288
rect 3700 8236 3752 8288
rect 4988 8236 5040 8288
rect 11336 8236 11388 8288
rect 11980 8236 12032 8288
rect 15108 8236 15160 8288
rect 15200 8236 15252 8288
rect 15844 8236 15896 8288
rect 17776 8304 17828 8356
rect 18972 8236 19024 8288
rect 3169 8134 3221 8186
rect 3233 8134 3285 8186
rect 3297 8134 3349 8186
rect 3361 8134 3413 8186
rect 3425 8134 3477 8186
rect 7608 8134 7660 8186
rect 7672 8134 7724 8186
rect 7736 8134 7788 8186
rect 7800 8134 7852 8186
rect 7864 8134 7916 8186
rect 12047 8134 12099 8186
rect 12111 8134 12163 8186
rect 12175 8134 12227 8186
rect 12239 8134 12291 8186
rect 12303 8134 12355 8186
rect 16486 8134 16538 8186
rect 16550 8134 16602 8186
rect 16614 8134 16666 8186
rect 16678 8134 16730 8186
rect 16742 8134 16794 8186
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 848 7828 900 7880
rect 1768 7828 1820 7880
rect 2136 7964 2188 8016
rect 2596 7964 2648 8016
rect 2320 7896 2372 7948
rect 6184 8032 6236 8084
rect 6368 8075 6420 8084
rect 6368 8041 6377 8075
rect 6377 8041 6411 8075
rect 6411 8041 6420 8075
rect 6368 8032 6420 8041
rect 7104 8032 7156 8084
rect 8576 8032 8628 8084
rect 3608 7828 3660 7880
rect 4344 7828 4396 7880
rect 12072 8032 12124 8084
rect 12256 8032 12308 8084
rect 12532 8032 12584 8084
rect 13452 8032 13504 8084
rect 13820 8032 13872 8084
rect 14372 8032 14424 8084
rect 15752 8032 15804 8084
rect 16028 8032 16080 8084
rect 16396 8032 16448 8084
rect 17040 8032 17092 8084
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 2136 7803 2188 7812
rect 2136 7769 2145 7803
rect 2145 7769 2179 7803
rect 2179 7769 2188 7803
rect 2136 7760 2188 7769
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 8392 7828 8444 7880
rect 9404 7896 9456 7948
rect 9496 7939 9548 7948
rect 9496 7905 9505 7939
rect 9505 7905 9539 7939
rect 9539 7905 9548 7939
rect 9496 7896 9548 7905
rect 11336 7964 11388 8016
rect 9864 7896 9916 7948
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 1308 7692 1360 7744
rect 5448 7760 5500 7812
rect 6000 7760 6052 7812
rect 4344 7692 4396 7744
rect 5908 7735 5960 7744
rect 5908 7701 5917 7735
rect 5917 7701 5951 7735
rect 5951 7701 5960 7735
rect 5908 7692 5960 7701
rect 6828 7692 6880 7744
rect 9036 7692 9088 7744
rect 10416 7760 10468 7812
rect 11152 7828 11204 7880
rect 11980 7828 12032 7880
rect 12716 7760 12768 7812
rect 9772 7692 9824 7744
rect 9956 7692 10008 7744
rect 10232 7692 10284 7744
rect 10508 7692 10560 7744
rect 10876 7692 10928 7744
rect 11336 7735 11388 7744
rect 11336 7701 11345 7735
rect 11345 7701 11379 7735
rect 11379 7701 11388 7735
rect 11336 7692 11388 7701
rect 11520 7692 11572 7744
rect 11612 7735 11664 7744
rect 11612 7701 11621 7735
rect 11621 7701 11655 7735
rect 11655 7701 11664 7735
rect 11612 7692 11664 7701
rect 12256 7692 12308 7744
rect 12808 7692 12860 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 13728 7896 13780 7948
rect 15016 8007 15068 8016
rect 15016 7973 15025 8007
rect 15025 7973 15059 8007
rect 15059 7973 15068 8007
rect 15016 7964 15068 7973
rect 17316 7964 17368 8016
rect 18420 7964 18472 8016
rect 15568 7896 15620 7948
rect 14740 7828 14792 7880
rect 14924 7760 14976 7812
rect 15108 7760 15160 7812
rect 15568 7760 15620 7812
rect 16856 7760 16908 7812
rect 17500 7828 17552 7880
rect 14096 7692 14148 7744
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 17132 7735 17184 7744
rect 17132 7701 17141 7735
rect 17141 7701 17175 7735
rect 17175 7701 17184 7735
rect 17132 7692 17184 7701
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 18236 7692 18288 7744
rect 3829 7590 3881 7642
rect 3893 7590 3945 7642
rect 3957 7590 4009 7642
rect 4021 7590 4073 7642
rect 4085 7590 4137 7642
rect 8268 7590 8320 7642
rect 8332 7590 8384 7642
rect 8396 7590 8448 7642
rect 8460 7590 8512 7642
rect 8524 7590 8576 7642
rect 12707 7590 12759 7642
rect 12771 7590 12823 7642
rect 12835 7590 12887 7642
rect 12899 7590 12951 7642
rect 12963 7590 13015 7642
rect 17146 7590 17198 7642
rect 17210 7590 17262 7642
rect 17274 7590 17326 7642
rect 17338 7590 17390 7642
rect 17402 7590 17454 7642
rect 388 7488 440 7540
rect 3424 7420 3476 7472
rect 3700 7488 3752 7540
rect 9772 7488 9824 7540
rect 9956 7488 10008 7540
rect 5816 7420 5868 7472
rect 9588 7463 9640 7472
rect 9588 7429 9597 7463
rect 9597 7429 9631 7463
rect 9631 7429 9640 7463
rect 9588 7420 9640 7429
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 5080 7352 5132 7404
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 1768 7284 1820 7336
rect 3516 7148 3568 7200
rect 9588 7284 9640 7336
rect 10508 7420 10560 7472
rect 12624 7488 12676 7540
rect 14188 7488 14240 7540
rect 14372 7531 14424 7540
rect 14372 7497 14381 7531
rect 14381 7497 14415 7531
rect 14415 7497 14424 7531
rect 14372 7488 14424 7497
rect 15476 7488 15528 7540
rect 15844 7488 15896 7540
rect 16028 7488 16080 7540
rect 17040 7488 17092 7540
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 18236 7488 18288 7540
rect 19248 7488 19300 7540
rect 15752 7420 15804 7472
rect 10600 7385 10609 7404
rect 10609 7385 10643 7404
rect 10643 7385 10652 7404
rect 10600 7352 10652 7385
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 12164 7395 12216 7404
rect 12164 7361 12173 7395
rect 12173 7361 12207 7395
rect 12207 7361 12216 7395
rect 12164 7352 12216 7361
rect 13452 7352 13504 7404
rect 15016 7352 15068 7404
rect 16304 7420 16356 7472
rect 17960 7420 18012 7472
rect 17132 7352 17184 7404
rect 18420 7352 18472 7404
rect 13176 7284 13228 7336
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 16028 7327 16080 7336
rect 16028 7293 16037 7327
rect 16037 7293 16071 7327
rect 16071 7293 16080 7327
rect 16028 7284 16080 7293
rect 17316 7284 17368 7336
rect 17408 7284 17460 7336
rect 4804 7216 4856 7268
rect 8300 7216 8352 7268
rect 9956 7216 10008 7268
rect 9772 7148 9824 7200
rect 11520 7216 11572 7268
rect 11980 7216 12032 7268
rect 12072 7216 12124 7268
rect 12900 7216 12952 7268
rect 13544 7216 13596 7268
rect 13728 7216 13780 7268
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 18788 7284 18840 7336
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 2320 6944 2372 6996
rect 6920 6944 6972 6996
rect 10508 6944 10560 6996
rect 11704 6944 11756 6996
rect 12164 6944 12216 6996
rect 12992 6944 13044 6996
rect 13360 6944 13412 6996
rect 15568 6944 15620 6996
rect 16304 6944 16356 6996
rect 17316 6944 17368 6996
rect 1768 6876 1820 6928
rect 2688 6876 2740 6928
rect 1400 6808 1452 6860
rect 8300 6876 8352 6928
rect 12716 6919 12768 6928
rect 12716 6885 12725 6919
rect 12725 6885 12759 6919
rect 12759 6885 12768 6919
rect 12716 6876 12768 6885
rect 12900 6876 12952 6928
rect 13728 6876 13780 6928
rect 15936 6876 15988 6928
rect 1860 6783 1912 6792
rect 1860 6749 1869 6783
rect 1869 6749 1903 6783
rect 1903 6749 1912 6783
rect 1860 6740 1912 6749
rect 2320 6740 2372 6792
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 2964 6740 3016 6792
rect 6736 6808 6788 6860
rect 9312 6808 9364 6860
rect 13636 6808 13688 6860
rect 16396 6808 16448 6860
rect 17592 6808 17644 6860
rect 2136 6715 2188 6724
rect 2136 6681 2145 6715
rect 2145 6681 2179 6715
rect 2179 6681 2188 6715
rect 2136 6672 2188 6681
rect 2504 6672 2556 6724
rect 1676 6647 1728 6656
rect 1676 6613 1685 6647
rect 1685 6613 1719 6647
rect 1719 6613 1728 6647
rect 1676 6604 1728 6613
rect 2780 6604 2832 6656
rect 2964 6647 3016 6656
rect 2964 6613 2973 6647
rect 2973 6613 3007 6647
rect 3007 6613 3016 6647
rect 2964 6604 3016 6613
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 3608 6672 3660 6724
rect 4068 6715 4120 6724
rect 4068 6681 4077 6715
rect 4077 6681 4111 6715
rect 4111 6681 4120 6715
rect 4068 6672 4120 6681
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 5632 6672 5684 6724
rect 7196 6672 7248 6724
rect 8668 6740 8720 6792
rect 10784 6740 10836 6792
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 12532 6740 12584 6792
rect 3700 6604 3752 6656
rect 9588 6604 9640 6656
rect 11796 6672 11848 6724
rect 12164 6672 12216 6724
rect 12256 6715 12308 6724
rect 12256 6681 12265 6715
rect 12265 6681 12299 6715
rect 12299 6681 12308 6715
rect 12256 6672 12308 6681
rect 12348 6672 12400 6724
rect 12992 6740 13044 6792
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 14096 6740 14148 6792
rect 17684 6740 17736 6792
rect 18052 6740 18104 6792
rect 11060 6604 11112 6656
rect 11244 6604 11296 6656
rect 12716 6604 12768 6656
rect 16856 6672 16908 6724
rect 17316 6672 17368 6724
rect 13820 6604 13872 6656
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 3829 6502 3881 6554
rect 3893 6502 3945 6554
rect 3957 6502 4009 6554
rect 4021 6502 4073 6554
rect 4085 6502 4137 6554
rect 8268 6502 8320 6554
rect 8332 6502 8384 6554
rect 8396 6502 8448 6554
rect 8460 6502 8512 6554
rect 8524 6502 8576 6554
rect 12707 6502 12759 6554
rect 12771 6502 12823 6554
rect 12835 6502 12887 6554
rect 12899 6502 12951 6554
rect 12963 6502 13015 6554
rect 17146 6502 17198 6554
rect 17210 6502 17262 6554
rect 17274 6502 17326 6554
rect 17338 6502 17390 6554
rect 17402 6502 17454 6554
rect 5172 6400 5224 6452
rect 1124 6332 1176 6384
rect 1400 6264 1452 6316
rect 2320 6332 2372 6384
rect 4528 6332 4580 6384
rect 4160 6264 4212 6316
rect 848 6196 900 6248
rect 2872 6128 2924 6180
rect 3700 6171 3752 6180
rect 3700 6137 3709 6171
rect 3709 6137 3743 6171
rect 3743 6137 3752 6171
rect 3700 6128 3752 6137
rect 1860 6060 1912 6112
rect 2964 6060 3016 6112
rect 4252 6196 4304 6248
rect 5632 6375 5684 6384
rect 5632 6341 5641 6375
rect 5641 6341 5675 6375
rect 5675 6341 5684 6375
rect 5632 6332 5684 6341
rect 5172 6264 5224 6316
rect 6552 6400 6604 6452
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 6736 6443 6788 6452
rect 6736 6409 6745 6443
rect 6745 6409 6779 6443
rect 6779 6409 6788 6443
rect 6736 6400 6788 6409
rect 7104 6443 7156 6452
rect 7104 6409 7113 6443
rect 7113 6409 7147 6443
rect 7147 6409 7156 6443
rect 7104 6400 7156 6409
rect 8392 6400 8444 6452
rect 9312 6400 9364 6452
rect 9404 6400 9456 6452
rect 10140 6400 10192 6452
rect 11244 6400 11296 6452
rect 11428 6400 11480 6452
rect 5816 6196 5868 6248
rect 4344 6128 4396 6180
rect 4896 6128 4948 6180
rect 6000 6128 6052 6180
rect 8116 6332 8168 6384
rect 9128 6375 9180 6384
rect 9128 6341 9137 6375
rect 9137 6341 9171 6375
rect 9171 6341 9180 6375
rect 9128 6332 9180 6341
rect 9496 6375 9548 6384
rect 9496 6341 9505 6375
rect 9505 6341 9539 6375
rect 9539 6341 9548 6375
rect 9496 6332 9548 6341
rect 10048 6375 10100 6384
rect 10048 6341 10057 6375
rect 10057 6341 10091 6375
rect 10091 6341 10100 6375
rect 10048 6332 10100 6341
rect 13084 6400 13136 6452
rect 14740 6400 14792 6452
rect 17040 6443 17092 6452
rect 17040 6409 17049 6443
rect 17049 6409 17083 6443
rect 17083 6409 17092 6443
rect 17040 6400 17092 6409
rect 17776 6400 17828 6452
rect 18512 6400 18564 6452
rect 9772 6264 9824 6316
rect 10600 6264 10652 6316
rect 11520 6264 11572 6316
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 7472 6196 7524 6248
rect 8760 6196 8812 6248
rect 12624 6332 12676 6384
rect 11888 6264 11940 6316
rect 12532 6307 12584 6316
rect 12532 6273 12541 6307
rect 12541 6273 12575 6307
rect 12575 6273 12584 6307
rect 12532 6264 12584 6273
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 12992 6196 13044 6248
rect 14004 6264 14056 6316
rect 6920 6128 6972 6180
rect 6828 6060 6880 6112
rect 7656 6171 7708 6180
rect 7656 6137 7665 6171
rect 7665 6137 7699 6171
rect 7699 6137 7708 6171
rect 7656 6128 7708 6137
rect 8116 6128 8168 6180
rect 10140 6128 10192 6180
rect 12072 6128 12124 6180
rect 16028 6128 16080 6180
rect 18420 6060 18472 6112
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 2228 5856 2280 5908
rect 2504 5856 2556 5908
rect 2872 5856 2924 5908
rect 4712 5856 4764 5908
rect 6000 5856 6052 5908
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 6460 5856 6512 5908
rect 2044 5788 2096 5840
rect 2412 5720 2464 5772
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2320 5652 2372 5704
rect 5540 5652 5592 5704
rect 6000 5652 6052 5704
rect 6368 5720 6420 5772
rect 8392 5856 8444 5908
rect 12532 5856 12584 5908
rect 13544 5856 13596 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 8484 5788 8536 5840
rect 10324 5788 10376 5840
rect 11152 5788 11204 5840
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 4160 5584 4212 5636
rect 5172 5584 5224 5636
rect 6460 5584 6512 5636
rect 8576 5720 8628 5772
rect 10232 5720 10284 5772
rect 10692 5720 10744 5772
rect 9956 5652 10008 5704
rect 11888 5652 11940 5704
rect 12624 5788 12676 5840
rect 16856 5856 16908 5908
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 18420 5856 18472 5908
rect 18880 5856 18932 5908
rect 12808 5720 12860 5772
rect 13084 5720 13136 5772
rect 13636 5720 13688 5772
rect 18052 5720 18104 5772
rect 14004 5652 14056 5704
rect 8024 5584 8076 5636
rect 8484 5584 8536 5636
rect 9404 5627 9456 5636
rect 9404 5593 9413 5627
rect 9413 5593 9447 5627
rect 9447 5593 9456 5627
rect 9404 5584 9456 5593
rect 2872 5516 2924 5568
rect 5080 5516 5132 5568
rect 5908 5516 5960 5568
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 10600 5584 10652 5636
rect 11244 5584 11296 5636
rect 14096 5584 14148 5636
rect 15108 5584 15160 5636
rect 7472 5516 7524 5525
rect 11704 5516 11756 5568
rect 12992 5516 13044 5568
rect 13912 5516 13964 5568
rect 3829 5414 3881 5466
rect 3893 5414 3945 5466
rect 3957 5414 4009 5466
rect 4021 5414 4073 5466
rect 4085 5414 4137 5466
rect 8268 5414 8320 5466
rect 8332 5414 8384 5466
rect 8396 5414 8448 5466
rect 8460 5414 8512 5466
rect 8524 5414 8576 5466
rect 12707 5414 12759 5466
rect 12771 5414 12823 5466
rect 12835 5414 12887 5466
rect 12899 5414 12951 5466
rect 12963 5414 13015 5466
rect 17146 5414 17198 5466
rect 17210 5414 17262 5466
rect 17274 5414 17326 5466
rect 17338 5414 17390 5466
rect 17402 5414 17454 5466
rect 2320 5355 2372 5364
rect 2320 5321 2329 5355
rect 2329 5321 2363 5355
rect 2363 5321 2372 5355
rect 2320 5312 2372 5321
rect 2596 5176 2648 5228
rect 2872 5176 2924 5228
rect 2964 5219 3016 5228
rect 2964 5185 2973 5219
rect 2973 5185 3007 5219
rect 3007 5185 3016 5219
rect 2964 5176 3016 5185
rect 848 5108 900 5160
rect 4160 5312 4212 5364
rect 4252 5312 4304 5364
rect 9220 5312 9272 5364
rect 9404 5312 9456 5364
rect 17960 5312 18012 5364
rect 4804 5244 4856 5296
rect 7012 5244 7064 5296
rect 15660 5244 15712 5296
rect 5724 5176 5776 5228
rect 6736 5176 6788 5228
rect 6644 5108 6696 5160
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 3516 4972 3568 5024
rect 4160 4972 4212 5024
rect 5356 5040 5408 5092
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 6368 4972 6420 5024
rect 6552 4972 6604 5024
rect 8024 5151 8076 5160
rect 8024 5117 8033 5151
rect 8033 5117 8067 5151
rect 8067 5117 8076 5151
rect 8024 5108 8076 5117
rect 8484 5108 8536 5160
rect 18696 5244 18748 5296
rect 18328 5219 18380 5228
rect 18328 5185 18337 5219
rect 18337 5185 18371 5219
rect 18371 5185 18380 5219
rect 18328 5176 18380 5185
rect 18420 5219 18472 5228
rect 18420 5185 18429 5219
rect 18429 5185 18463 5219
rect 18463 5185 18472 5219
rect 18420 5176 18472 5185
rect 16304 5108 16356 5160
rect 17868 5040 17920 5092
rect 14832 4972 14884 5024
rect 18052 4972 18104 5024
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 2044 4768 2096 4820
rect 2596 4811 2648 4820
rect 2596 4777 2605 4811
rect 2605 4777 2639 4811
rect 2639 4777 2648 4811
rect 2596 4768 2648 4777
rect 2964 4768 3016 4820
rect 4160 4768 4212 4820
rect 4988 4768 5040 4820
rect 2872 4700 2924 4752
rect 3884 4700 3936 4752
rect 6460 4700 6512 4752
rect 6644 4700 6696 4752
rect 8484 4700 8536 4752
rect 13176 4768 13228 4820
rect 7288 4632 7340 4684
rect 9680 4632 9732 4684
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4344 4564 4396 4616
rect 4804 4564 4856 4616
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 14372 4700 14424 4752
rect 14096 4632 14148 4684
rect 14832 4768 14884 4820
rect 19156 4700 19208 4752
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 14464 4564 14516 4616
rect 848 4496 900 4548
rect 3332 4496 3384 4548
rect 13084 4496 13136 4548
rect 13636 4496 13688 4548
rect 16120 4496 16172 4548
rect 18144 4564 18196 4616
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 5264 4428 5316 4480
rect 17500 4428 17552 4480
rect 3829 4326 3881 4378
rect 3893 4326 3945 4378
rect 3957 4326 4009 4378
rect 4021 4326 4073 4378
rect 4085 4326 4137 4378
rect 8268 4326 8320 4378
rect 8332 4326 8384 4378
rect 8396 4326 8448 4378
rect 8460 4326 8512 4378
rect 8524 4326 8576 4378
rect 12707 4326 12759 4378
rect 12771 4326 12823 4378
rect 12835 4326 12887 4378
rect 12899 4326 12951 4378
rect 12963 4326 13015 4378
rect 17146 4326 17198 4378
rect 17210 4326 17262 4378
rect 17274 4326 17326 4378
rect 17338 4326 17390 4378
rect 17402 4326 17454 4378
rect 1860 4224 1912 4276
rect 3332 4224 3384 4276
rect 4344 4224 4396 4276
rect 4436 4224 4488 4276
rect 8852 4224 8904 4276
rect 9772 4224 9824 4276
rect 2780 4088 2832 4140
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 5540 4156 5592 4208
rect 10784 4156 10836 4208
rect 13820 4224 13872 4276
rect 4436 4063 4488 4072
rect 4436 4029 4445 4063
rect 4445 4029 4479 4063
rect 4479 4029 4488 4063
rect 4436 4020 4488 4029
rect 6276 4088 6328 4140
rect 7472 4088 7524 4140
rect 8944 4088 8996 4140
rect 15108 4156 15160 4208
rect 17408 4156 17460 4208
rect 13084 4088 13136 4140
rect 756 3952 808 4004
rect 3516 3884 3568 3936
rect 6184 3952 6236 4004
rect 9036 3952 9088 4004
rect 12624 4020 12676 4072
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 11152 3884 11204 3936
rect 11612 3884 11664 3936
rect 13360 3884 13412 3936
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 15476 4088 15528 4140
rect 16396 4088 16448 4140
rect 17868 4088 17920 4140
rect 14280 4020 14332 4072
rect 16304 4020 16356 4072
rect 16396 3927 16448 3936
rect 16396 3893 16405 3927
rect 16405 3893 16439 3927
rect 16439 3893 16448 3927
rect 16396 3884 16448 3893
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 2964 3723 3016 3732
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 3700 3612 3752 3664
rect 4436 3680 4488 3732
rect 5724 3680 5776 3732
rect 6460 3723 6512 3732
rect 6460 3689 6469 3723
rect 6469 3689 6503 3723
rect 6503 3689 6512 3723
rect 6460 3680 6512 3689
rect 10048 3680 10100 3732
rect 10416 3680 10468 3732
rect 11152 3680 11204 3732
rect 11336 3680 11388 3732
rect 8760 3612 8812 3664
rect 12348 3612 12400 3664
rect 848 3544 900 3596
rect 2964 3544 3016 3596
rect 11796 3544 11848 3596
rect 13636 3723 13688 3732
rect 13636 3689 13645 3723
rect 13645 3689 13679 3723
rect 13679 3689 13688 3723
rect 13636 3680 13688 3689
rect 13176 3612 13228 3664
rect 15016 3680 15068 3732
rect 15200 3723 15252 3732
rect 15200 3689 15209 3723
rect 15209 3689 15243 3723
rect 15243 3689 15252 3723
rect 15200 3680 15252 3689
rect 15476 3723 15528 3732
rect 15476 3689 15485 3723
rect 15485 3689 15519 3723
rect 15519 3689 15528 3723
rect 15476 3680 15528 3689
rect 14648 3655 14700 3664
rect 14648 3621 14657 3655
rect 14657 3621 14691 3655
rect 14691 3621 14700 3655
rect 14648 3612 14700 3621
rect 3056 3476 3108 3528
rect 5540 3519 5592 3528
rect 5540 3485 5548 3519
rect 5548 3485 5582 3519
rect 5582 3485 5592 3519
rect 5540 3476 5592 3485
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 8668 3476 8720 3528
rect 10692 3476 10744 3528
rect 12624 3476 12676 3528
rect 13360 3544 13412 3596
rect 13728 3544 13780 3596
rect 14464 3544 14516 3596
rect 15844 3544 15896 3596
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 6092 3451 6144 3460
rect 6092 3417 6101 3451
rect 6101 3417 6135 3451
rect 6135 3417 6144 3451
rect 6092 3408 6144 3417
rect 6276 3408 6328 3460
rect 10048 3408 10100 3460
rect 10784 3408 10836 3460
rect 11152 3408 11204 3460
rect 2136 3383 2188 3392
rect 2136 3349 2145 3383
rect 2145 3349 2179 3383
rect 2179 3349 2188 3383
rect 2136 3340 2188 3349
rect 2504 3340 2556 3392
rect 4436 3340 4488 3392
rect 4528 3340 4580 3392
rect 5356 3340 5408 3392
rect 7840 3383 7892 3392
rect 7840 3349 7849 3383
rect 7849 3349 7883 3383
rect 7883 3349 7892 3383
rect 7840 3340 7892 3349
rect 8668 3340 8720 3392
rect 9036 3340 9088 3392
rect 12348 3340 12400 3392
rect 14096 3408 14148 3460
rect 16212 3476 16264 3528
rect 15568 3408 15620 3460
rect 15936 3383 15988 3392
rect 15936 3349 15945 3383
rect 15945 3349 15979 3383
rect 15979 3349 15988 3383
rect 15936 3340 15988 3349
rect 16396 3340 16448 3392
rect 17408 3340 17460 3392
rect 3829 3238 3881 3290
rect 3893 3238 3945 3290
rect 3957 3238 4009 3290
rect 4021 3238 4073 3290
rect 4085 3238 4137 3290
rect 8268 3238 8320 3290
rect 8332 3238 8384 3290
rect 8396 3238 8448 3290
rect 8460 3238 8512 3290
rect 8524 3238 8576 3290
rect 12707 3238 12759 3290
rect 12771 3238 12823 3290
rect 12835 3238 12887 3290
rect 12899 3238 12951 3290
rect 12963 3238 13015 3290
rect 17146 3238 17198 3290
rect 17210 3238 17262 3290
rect 17274 3238 17326 3290
rect 17338 3238 17390 3290
rect 17402 3238 17454 3290
rect 1768 3136 1820 3188
rect 3148 3136 3200 3188
rect 3608 3136 3660 3188
rect 4528 3136 4580 3188
rect 4896 3136 4948 3188
rect 5356 3136 5408 3188
rect 5540 3136 5592 3188
rect 6000 3136 6052 3188
rect 7472 3179 7524 3188
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 10324 3179 10376 3188
rect 10324 3145 10333 3179
rect 10333 3145 10367 3179
rect 10367 3145 10376 3179
rect 10324 3136 10376 3145
rect 12532 3179 12584 3188
rect 12532 3145 12541 3179
rect 12541 3145 12575 3179
rect 12575 3145 12584 3179
rect 12532 3136 12584 3145
rect 12624 3136 12676 3188
rect 13360 3136 13412 3188
rect 15292 3136 15344 3188
rect 15844 3136 15896 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 2688 3000 2740 3052
rect 848 2932 900 2984
rect 3148 2864 3200 2916
rect 7932 3068 7984 3120
rect 5448 3000 5500 3052
rect 6276 2932 6328 2984
rect 7380 2932 7432 2984
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 8760 3000 8812 3052
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 9588 3000 9640 3052
rect 14924 3068 14976 3120
rect 16396 3068 16448 3120
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 8300 2932 8352 2984
rect 9680 2932 9732 2984
rect 10324 2932 10376 2984
rect 9864 2864 9916 2916
rect 10140 2864 10192 2916
rect 11612 2932 11664 2984
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 13176 3000 13228 3052
rect 12624 2932 12676 2984
rect 13084 2932 13136 2984
rect 13452 2932 13504 2984
rect 14096 2932 14148 2984
rect 17408 2932 17460 2984
rect 18420 3000 18472 3052
rect 19340 2932 19392 2984
rect 6828 2796 6880 2848
rect 8760 2796 8812 2848
rect 11060 2796 11112 2848
rect 15936 2864 15988 2916
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 1492 2592 1544 2644
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 6552 2592 6604 2644
rect 940 2524 992 2576
rect 7196 2524 7248 2576
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 10232 2592 10284 2644
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 11152 2592 11204 2644
rect 8760 2567 8812 2576
rect 8760 2533 8769 2567
rect 8769 2533 8803 2567
rect 8803 2533 8812 2567
rect 8760 2524 8812 2533
rect 8944 2524 8996 2576
rect 13360 2592 13412 2644
rect 14004 2592 14056 2644
rect 14372 2592 14424 2644
rect 17316 2635 17368 2644
rect 17316 2601 17325 2635
rect 17325 2601 17359 2635
rect 17359 2601 17368 2635
rect 17316 2592 17368 2601
rect 18604 2592 18656 2644
rect 14464 2524 14516 2576
rect 14924 2524 14976 2576
rect 8300 2456 8352 2508
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 2872 2431 2924 2440
rect 848 2320 900 2372
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 4804 2388 4856 2440
rect 7748 2388 7800 2440
rect 8668 2388 8720 2440
rect 9036 2388 9088 2440
rect 9680 2388 9732 2440
rect 2780 2320 2832 2372
rect 5264 2252 5316 2304
rect 9220 2252 9272 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 12624 2456 12676 2508
rect 12808 2456 12860 2508
rect 10324 2388 10376 2440
rect 11060 2388 11112 2440
rect 12072 2363 12124 2372
rect 12072 2329 12081 2363
rect 12081 2329 12115 2363
rect 12115 2329 12124 2363
rect 12072 2320 12124 2329
rect 13820 2320 13872 2372
rect 12808 2252 12860 2304
rect 13360 2252 13412 2304
rect 14556 2388 14608 2440
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 18236 2524 18288 2576
rect 19432 2388 19484 2440
rect 18788 2320 18840 2372
rect 3829 2150 3881 2202
rect 3893 2150 3945 2202
rect 3957 2150 4009 2202
rect 4021 2150 4073 2202
rect 4085 2150 4137 2202
rect 8268 2150 8320 2202
rect 8332 2150 8384 2202
rect 8396 2150 8448 2202
rect 8460 2150 8512 2202
rect 8524 2150 8576 2202
rect 12707 2150 12759 2202
rect 12771 2150 12823 2202
rect 12835 2150 12887 2202
rect 12899 2150 12951 2202
rect 12963 2150 13015 2202
rect 17146 2150 17198 2202
rect 17210 2150 17262 2202
rect 17274 2150 17326 2202
rect 17338 2150 17390 2202
rect 17402 2150 17454 2202
rect 8116 2048 8168 2100
rect 15108 2048 15160 2100
rect 9220 1980 9272 2032
rect 11704 1980 11756 2032
rect 7196 1912 7248 1964
rect 11244 1912 11296 1964
rect 572 1844 624 1896
rect 12072 1844 12124 1896
<< metal2 >>
rect 2870 19136 2926 19145
rect 2870 19071 2926 19080
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 938 17912 994 17921
rect 938 17847 994 17856
rect 952 16697 980 17847
rect 2792 17354 2820 18391
rect 2700 17326 2820 17354
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 386 16688 442 16697
rect 386 16623 442 16632
rect 938 16688 994 16697
rect 938 16623 994 16632
rect 400 7546 428 16623
rect 1504 16425 1532 17138
rect 2700 17134 2728 17326
rect 2884 17270 2912 19071
rect 6734 18184 6790 18193
rect 6734 18119 6790 18128
rect 2962 17776 3018 17785
rect 2962 17711 3018 17720
rect 2976 17270 3004 17711
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 3829 17436 4137 17445
rect 3829 17434 3835 17436
rect 3891 17434 3915 17436
rect 3971 17434 3995 17436
rect 4051 17434 4075 17436
rect 4131 17434 4137 17436
rect 3891 17382 3893 17434
rect 4073 17382 4075 17434
rect 3829 17380 3835 17382
rect 3891 17380 3915 17382
rect 3971 17380 3995 17382
rect 4051 17380 4075 17382
rect 4131 17380 4137 17382
rect 3829 17371 4137 17380
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 3608 17264 3660 17270
rect 3608 17206 3660 17212
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1964 16590 1992 17002
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1860 16448 1912 16454
rect 1490 16416 1546 16425
rect 1860 16390 1912 16396
rect 1490 16351 1546 16360
rect 848 16040 900 16046
rect 848 15982 900 15988
rect 860 15881 888 15982
rect 846 15872 902 15881
rect 846 15807 902 15816
rect 1504 15502 1532 16351
rect 1676 15564 1728 15570
rect 1676 15506 1728 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1492 15496 1544 15502
rect 1492 15438 1544 15444
rect 940 15360 992 15366
rect 940 15302 992 15308
rect 756 14340 808 14346
rect 756 14282 808 14288
rect 572 11892 624 11898
rect 572 11834 624 11840
rect 388 7540 440 7546
rect 388 7482 440 7488
rect 584 1902 612 11834
rect 768 4010 796 14282
rect 848 12300 900 12306
rect 848 12242 900 12248
rect 860 7886 888 12242
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 848 6248 900 6254
rect 848 6190 900 6196
rect 860 6089 888 6190
rect 846 6080 902 6089
rect 846 6015 902 6024
rect 848 5160 900 5166
rect 848 5102 900 5108
rect 860 5001 888 5102
rect 846 4992 902 5001
rect 846 4927 902 4936
rect 848 4548 900 4554
rect 848 4490 900 4496
rect 860 4321 888 4490
rect 846 4312 902 4321
rect 846 4247 902 4256
rect 756 4004 808 4010
rect 756 3946 808 3952
rect 846 3632 902 3641
rect 846 3567 848 3576
rect 900 3567 902 3576
rect 848 3538 900 3544
rect 848 2984 900 2990
rect 846 2952 848 2961
rect 900 2952 902 2961
rect 846 2887 902 2896
rect 952 2582 980 15302
rect 1412 15065 1440 15438
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1492 15020 1544 15026
rect 1412 14618 1440 14991
rect 1492 14962 1544 14968
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1504 14482 1532 14962
rect 1688 14958 1716 15506
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1216 14408 1268 14414
rect 1214 14376 1216 14385
rect 1268 14376 1270 14385
rect 1214 14311 1270 14320
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1214 12880 1270 12889
rect 1214 12815 1270 12824
rect 1032 12640 1084 12646
rect 1032 12582 1084 12588
rect 1044 4729 1072 12582
rect 1228 12306 1256 12815
rect 1412 12345 1440 13262
rect 1398 12336 1454 12345
rect 1216 12300 1268 12306
rect 1398 12271 1454 12280
rect 1504 12322 1532 14418
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1596 14278 1624 14311
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1596 13977 1624 14010
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 1688 13326 1716 14214
rect 1872 13326 1900 16390
rect 1964 14550 1992 16526
rect 2056 14890 2084 16594
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 2134 16008 2190 16017
rect 2134 15943 2190 15952
rect 2044 14884 2096 14890
rect 2044 14826 2096 14832
rect 1952 14544 2004 14550
rect 1952 14486 2004 14492
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13326 1992 13670
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1582 12336 1638 12345
rect 1504 12294 1582 12322
rect 1216 12242 1268 12248
rect 1124 12232 1176 12238
rect 1124 12174 1176 12180
rect 1214 12200 1270 12209
rect 1136 6390 1164 12174
rect 1214 12135 1270 12144
rect 1228 8362 1256 12135
rect 1308 11280 1360 11286
rect 1308 11222 1360 11228
rect 1216 8356 1268 8362
rect 1216 8298 1268 8304
rect 1320 7750 1348 11222
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10305 1440 10610
rect 1398 10296 1454 10305
rect 1398 10231 1400 10240
rect 1452 10231 1454 10240
rect 1400 10202 1452 10208
rect 1504 9081 1532 12294
rect 1582 12271 1638 12280
rect 1584 12164 1636 12170
rect 1584 12106 1636 12112
rect 1596 11665 1624 12106
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11762 1716 12038
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1582 11656 1638 11665
rect 1582 11591 1638 11600
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 10742 1624 11494
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1584 10736 1636 10742
rect 1584 10678 1636 10684
rect 1582 10568 1638 10577
rect 1582 10503 1584 10512
rect 1636 10503 1638 10512
rect 1584 10474 1636 10480
rect 1688 10146 1716 11018
rect 1596 10118 1716 10146
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1400 8968 1452 8974
rect 1398 8936 1400 8945
rect 1452 8936 1454 8945
rect 1398 8871 1454 8880
rect 1596 8786 1624 10118
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1412 8758 1624 8786
rect 1308 7744 1360 7750
rect 1308 7686 1360 7692
rect 1412 6866 1440 8758
rect 1490 8664 1546 8673
rect 1490 8599 1546 8608
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1124 6384 1176 6390
rect 1124 6326 1176 6332
rect 1412 6322 1440 6802
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1030 4720 1086 4729
rect 1030 4655 1086 4664
rect 1504 2650 1532 8599
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1596 7954 1624 8191
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 6905 1624 7278
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1688 6746 1716 9998
rect 1780 9654 1808 13126
rect 1872 12782 1900 13126
rect 1964 13025 1992 13262
rect 1950 13016 2006 13025
rect 1950 12951 2006 12960
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1860 12368 1912 12374
rect 1860 12310 1912 12316
rect 1872 11558 1900 12310
rect 2056 12238 2084 13806
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 2056 11642 2084 12174
rect 2148 11762 2176 15943
rect 2240 14906 2268 16458
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2608 15570 2636 15982
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 2332 15162 2360 15370
rect 2412 15360 2464 15366
rect 2410 15328 2412 15337
rect 2464 15328 2466 15337
rect 2410 15263 2466 15272
rect 2700 15178 2728 16934
rect 2780 16584 2832 16590
rect 2778 16552 2780 16561
rect 2832 16552 2834 16561
rect 2778 16487 2834 16496
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 16153 2820 16390
rect 2778 16144 2834 16153
rect 2778 16079 2780 16088
rect 2832 16079 2834 16088
rect 2780 16050 2832 16056
rect 2884 15706 2912 17206
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3068 17105 3096 17138
rect 3516 17128 3568 17134
rect 3054 17096 3110 17105
rect 3516 17070 3568 17076
rect 3054 17031 3110 17040
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2976 16561 3004 16594
rect 2962 16552 3018 16561
rect 2962 16487 3018 16496
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2320 15156 2372 15162
rect 2700 15150 2912 15178
rect 2976 15162 3004 16050
rect 2320 15098 2372 15104
rect 2780 15088 2832 15094
rect 2502 15056 2558 15065
rect 2780 15030 2832 15036
rect 2502 14991 2558 15000
rect 2240 14878 2360 14906
rect 2226 14512 2282 14521
rect 2226 14447 2282 14456
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1964 11082 1992 11630
rect 2056 11614 2176 11642
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 10130 1900 10950
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1964 10198 1992 10678
rect 1952 10192 2004 10198
rect 1952 10134 2004 10140
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1872 9466 1900 10066
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1964 9625 1992 9998
rect 2056 9722 2084 11086
rect 2148 10690 2176 11614
rect 2240 10810 2268 14447
rect 2332 13190 2360 14878
rect 2412 14884 2464 14890
rect 2412 14826 2464 14832
rect 2424 13190 2452 14826
rect 2516 13530 2544 14991
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2700 14113 2728 14894
rect 2686 14104 2742 14113
rect 2686 14039 2742 14048
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2608 13274 2636 13670
rect 2516 13246 2636 13274
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2412 11756 2464 11762
rect 2516 11744 2544 13246
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 12306 2636 13126
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2464 11716 2544 11744
rect 2412 11698 2464 11704
rect 2318 11248 2374 11257
rect 2318 11183 2374 11192
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2148 10662 2268 10690
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2148 10198 2176 10542
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 1950 9616 2006 9625
rect 1950 9551 2006 9560
rect 1872 9438 1992 9466
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1780 7342 1808 7822
rect 1872 7449 1900 8230
rect 1858 7440 1914 7449
rect 1858 7375 1860 7384
rect 1912 7375 1914 7384
rect 1860 7346 1912 7352
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1780 6934 1808 7278
rect 1768 6928 1820 6934
rect 1768 6870 1820 6876
rect 1860 6792 1912 6798
rect 1688 6718 1808 6746
rect 1860 6734 1912 6740
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 5817 1716 6598
rect 1674 5808 1730 5817
rect 1674 5743 1730 5752
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1596 5545 1624 5578
rect 1582 5536 1638 5545
rect 1582 5471 1638 5480
rect 1780 3194 1808 6718
rect 1872 6118 1900 6734
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1964 5710 1992 9438
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 2056 5846 2084 8842
rect 2148 8022 2176 9998
rect 2240 9110 2268 10662
rect 2332 10470 2360 11183
rect 2424 10810 2452 11698
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2332 9178 2360 10406
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 9104 2280 9110
rect 2228 9046 2280 9052
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2148 7585 2176 7754
rect 2134 7576 2190 7585
rect 2134 7511 2190 7520
rect 2134 7304 2190 7313
rect 2134 7239 2190 7248
rect 2148 6730 2176 7239
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 2240 5914 2268 8910
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2332 7002 2360 7890
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2424 6905 2452 9930
rect 2516 8514 2544 11562
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2608 9178 2636 11154
rect 2700 11082 2728 12786
rect 2792 11762 2820 15030
rect 2884 13870 2912 15150
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2976 14482 3004 15098
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2884 12628 2912 13806
rect 2976 12986 3004 14418
rect 3068 13938 3096 16934
rect 3169 16892 3477 16901
rect 3169 16890 3175 16892
rect 3231 16890 3255 16892
rect 3311 16890 3335 16892
rect 3391 16890 3415 16892
rect 3471 16890 3477 16892
rect 3231 16838 3233 16890
rect 3413 16838 3415 16890
rect 3169 16836 3175 16838
rect 3231 16836 3255 16838
rect 3311 16836 3335 16838
rect 3391 16836 3415 16838
rect 3471 16836 3477 16838
rect 3169 16827 3477 16836
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3252 16046 3280 16594
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3169 15804 3477 15813
rect 3169 15802 3175 15804
rect 3231 15802 3255 15804
rect 3311 15802 3335 15804
rect 3391 15802 3415 15804
rect 3471 15802 3477 15804
rect 3231 15750 3233 15802
rect 3413 15750 3415 15802
rect 3169 15748 3175 15750
rect 3231 15748 3255 15750
rect 3311 15748 3335 15750
rect 3391 15748 3415 15750
rect 3471 15748 3477 15750
rect 3169 15739 3477 15748
rect 3528 15706 3556 17070
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3620 15502 3648 17206
rect 3712 16232 3740 17274
rect 4344 17264 4396 17270
rect 4396 17224 4476 17252
rect 4344 17206 4396 17212
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3804 16726 3832 16934
rect 3792 16720 3844 16726
rect 3896 16697 3924 16934
rect 4448 16794 4476 17224
rect 6012 17202 6040 17478
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5356 17128 5408 17134
rect 5078 17096 5134 17105
rect 5632 17128 5684 17134
rect 5408 17088 5580 17116
rect 5356 17070 5408 17076
rect 5078 17031 5134 17040
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4344 16720 4396 16726
rect 3792 16662 3844 16668
rect 3882 16688 3938 16697
rect 4344 16662 4396 16668
rect 3882 16623 3938 16632
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 3829 16348 4137 16357
rect 3829 16346 3835 16348
rect 3891 16346 3915 16348
rect 3971 16346 3995 16348
rect 4051 16346 4075 16348
rect 4131 16346 4137 16348
rect 3891 16294 3893 16346
rect 4073 16294 4075 16346
rect 3829 16292 3835 16294
rect 3891 16292 3915 16294
rect 3971 16292 3995 16294
rect 4051 16292 4075 16294
rect 4131 16292 4137 16294
rect 3829 16283 4137 16292
rect 3712 16204 3832 16232
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3148 15360 3200 15366
rect 3146 15328 3148 15337
rect 3200 15328 3202 15337
rect 3146 15263 3202 15272
rect 3344 14958 3372 15370
rect 3804 15348 3832 16204
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 3712 15320 3832 15348
rect 4080 15348 4108 16079
rect 4264 15434 4292 16594
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4080 15320 4200 15348
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3169 14716 3477 14725
rect 3169 14714 3175 14716
rect 3231 14714 3255 14716
rect 3311 14714 3335 14716
rect 3391 14714 3415 14716
rect 3471 14714 3477 14716
rect 3231 14662 3233 14714
rect 3413 14662 3415 14714
rect 3169 14660 3175 14662
rect 3231 14660 3255 14662
rect 3311 14660 3335 14662
rect 3391 14660 3415 14662
rect 3471 14660 3477 14662
rect 3169 14651 3477 14660
rect 3712 14006 3740 15320
rect 3829 15260 4137 15269
rect 3829 15258 3835 15260
rect 3891 15258 3915 15260
rect 3971 15258 3995 15260
rect 4051 15258 4075 15260
rect 4131 15258 4137 15260
rect 3891 15206 3893 15258
rect 4073 15206 4075 15258
rect 3829 15204 3835 15206
rect 3891 15204 3915 15206
rect 3971 15204 3995 15206
rect 4051 15204 4075 15206
rect 4131 15204 4137 15206
rect 3829 15195 4137 15204
rect 4172 15042 4200 15320
rect 4080 15014 4200 15042
rect 4080 14822 4108 15014
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4356 14362 4384 16662
rect 4448 16182 4476 16730
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4436 16176 4488 16182
rect 4436 16118 4488 16124
rect 4448 15094 4476 16118
rect 4632 15201 4660 16390
rect 4724 16114 4752 16526
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 5092 15706 5120 17031
rect 5552 16794 5580 17088
rect 5632 17070 5684 17076
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5262 16552 5318 16561
rect 5262 16487 5264 16496
rect 5316 16487 5318 16496
rect 5264 16458 5316 16464
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4618 15192 4674 15201
rect 4618 15127 4674 15136
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4436 14952 4488 14958
rect 4434 14920 4436 14929
rect 4488 14920 4490 14929
rect 4434 14855 4490 14864
rect 3976 14340 4028 14346
rect 4160 14340 4212 14346
rect 4028 14300 4160 14328
rect 3976 14282 4028 14288
rect 4160 14282 4212 14288
rect 4264 14334 4384 14362
rect 3829 14172 4137 14181
rect 3829 14170 3835 14172
rect 3891 14170 3915 14172
rect 3971 14170 3995 14172
rect 4051 14170 4075 14172
rect 4131 14170 4137 14172
rect 3891 14118 3893 14170
rect 4073 14118 4075 14170
rect 3829 14116 3835 14118
rect 3891 14116 3915 14118
rect 3971 14116 3995 14118
rect 4051 14116 4075 14118
rect 4131 14116 4137 14118
rect 3829 14107 4137 14116
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 13410 3096 13874
rect 3169 13628 3477 13637
rect 3169 13626 3175 13628
rect 3231 13626 3255 13628
rect 3311 13626 3335 13628
rect 3391 13626 3415 13628
rect 3471 13626 3477 13628
rect 3231 13574 3233 13626
rect 3413 13574 3415 13626
rect 3169 13572 3175 13574
rect 3231 13572 3255 13574
rect 3311 13572 3335 13574
rect 3391 13572 3415 13574
rect 3471 13572 3477 13574
rect 3169 13563 3477 13572
rect 3068 13382 3372 13410
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 3160 12730 3188 13262
rect 3068 12702 3188 12730
rect 2884 12600 3004 12628
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11830 2912 12038
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2700 9654 2728 9930
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2516 8486 2636 8514
rect 2608 8401 2636 8486
rect 2594 8392 2650 8401
rect 2594 8327 2650 8336
rect 2596 8016 2648 8022
rect 2700 7993 2728 9590
rect 2596 7958 2648 7964
rect 2686 7984 2742 7993
rect 2410 6896 2466 6905
rect 2410 6831 2466 6840
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2332 6390 2360 6734
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2318 6216 2374 6225
rect 2318 6151 2374 6160
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1872 4282 1900 4558
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1964 2774 1992 5646
rect 2056 4826 2084 5782
rect 2332 5710 2360 6151
rect 2424 5778 2452 6831
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2516 5914 2544 6666
rect 2608 6225 2636 7958
rect 2686 7919 2742 7928
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2594 6216 2650 6225
rect 2594 6151 2650 6160
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2332 5370 2360 5646
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2516 3398 2544 5850
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2608 5137 2636 5170
rect 2594 5128 2650 5137
rect 2594 5063 2650 5072
rect 2608 4826 2636 5063
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2148 3058 2176 3334
rect 2700 3058 2728 6870
rect 2792 6798 2820 11562
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2884 10470 2912 10610
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2884 9178 2912 10406
rect 2976 10130 3004 12600
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 4146 2820 6598
rect 2884 6186 2912 8978
rect 2976 8634 3004 10066
rect 3068 9994 3096 12702
rect 3344 12628 3372 13382
rect 3712 13326 3740 13942
rect 4160 13932 4212 13938
rect 4080 13892 4160 13920
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3988 13569 4016 13806
rect 3974 13560 4030 13569
rect 4080 13530 4108 13892
rect 4160 13874 4212 13880
rect 3974 13495 4030 13504
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 3700 13320 3752 13326
rect 3606 13288 3662 13297
rect 3700 13262 3752 13268
rect 3606 13223 3608 13232
rect 3660 13223 3662 13232
rect 3608 13194 3660 13200
rect 3829 13084 4137 13093
rect 3829 13082 3835 13084
rect 3891 13082 3915 13084
rect 3971 13082 3995 13084
rect 4051 13082 4075 13084
rect 4131 13082 4137 13084
rect 3891 13030 3893 13082
rect 4073 13030 4075 13082
rect 3829 13028 3835 13030
rect 3891 13028 3915 13030
rect 3971 13028 3995 13030
rect 4051 13028 4075 13030
rect 4131 13028 4137 13030
rect 3829 13019 4137 13028
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3436 12850 3464 12922
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3436 12730 3464 12786
rect 3436 12702 3648 12730
rect 3344 12600 3556 12628
rect 3169 12540 3477 12549
rect 3169 12538 3175 12540
rect 3231 12538 3255 12540
rect 3311 12538 3335 12540
rect 3391 12538 3415 12540
rect 3471 12538 3477 12540
rect 3231 12486 3233 12538
rect 3413 12486 3415 12538
rect 3169 12484 3175 12486
rect 3231 12484 3255 12486
rect 3311 12484 3335 12486
rect 3391 12484 3415 12486
rect 3471 12484 3477 12486
rect 3169 12475 3477 12484
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3160 11558 3188 12106
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3169 11452 3477 11461
rect 3169 11450 3175 11452
rect 3231 11450 3255 11452
rect 3311 11450 3335 11452
rect 3391 11450 3415 11452
rect 3471 11450 3477 11452
rect 3231 11398 3233 11450
rect 3413 11398 3415 11450
rect 3169 11396 3175 11398
rect 3231 11396 3255 11398
rect 3311 11396 3335 11398
rect 3391 11396 3415 11398
rect 3471 11396 3477 11398
rect 3169 11387 3477 11396
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3344 10713 3372 10746
rect 3330 10704 3386 10713
rect 3330 10639 3386 10648
rect 3436 10606 3464 10950
rect 3528 10724 3556 12600
rect 3620 12442 3648 12702
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3712 12481 3740 12582
rect 3698 12472 3754 12481
rect 3608 12436 3660 12442
rect 3698 12407 3754 12416
rect 3608 12378 3660 12384
rect 3804 12084 3832 12922
rect 4172 12646 4200 13330
rect 4264 13025 4292 14334
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4356 14113 4384 14214
rect 4342 14104 4398 14113
rect 4342 14039 4398 14048
rect 4356 13938 4384 14039
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4448 13818 4476 14855
rect 4356 13790 4476 13818
rect 4250 13016 4306 13025
rect 4250 12951 4306 12960
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3712 12056 3832 12084
rect 3712 11830 3740 12056
rect 3829 11996 4137 12005
rect 3829 11994 3835 11996
rect 3891 11994 3915 11996
rect 3971 11994 3995 11996
rect 4051 11994 4075 11996
rect 4131 11994 4137 11996
rect 3891 11942 3893 11994
rect 4073 11942 4075 11994
rect 3829 11940 3835 11942
rect 3891 11940 3915 11942
rect 3971 11940 3995 11942
rect 4051 11940 4075 11942
rect 4131 11940 4137 11942
rect 3829 11931 4137 11940
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3712 10792 3740 11766
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 11286 4016 11698
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4080 11014 4108 11766
rect 4172 11218 4200 12378
rect 4250 12336 4306 12345
rect 4250 12271 4306 12280
rect 4264 12238 4292 12271
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3829 10908 4137 10917
rect 3829 10906 3835 10908
rect 3891 10906 3915 10908
rect 3971 10906 3995 10908
rect 4051 10906 4075 10908
rect 4131 10906 4137 10908
rect 3891 10854 3893 10906
rect 4073 10854 4075 10906
rect 3829 10852 3835 10854
rect 3891 10852 3915 10854
rect 3971 10852 3995 10854
rect 4051 10852 4075 10854
rect 4131 10852 4137 10854
rect 3829 10843 4137 10852
rect 3712 10764 3832 10792
rect 3528 10696 3740 10724
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3169 10364 3477 10373
rect 3169 10362 3175 10364
rect 3231 10362 3255 10364
rect 3311 10362 3335 10364
rect 3391 10362 3415 10364
rect 3471 10362 3477 10364
rect 3231 10310 3233 10362
rect 3413 10310 3415 10362
rect 3169 10308 3175 10310
rect 3231 10308 3255 10310
rect 3311 10308 3335 10310
rect 3391 10308 3415 10310
rect 3471 10308 3477 10310
rect 3169 10299 3477 10308
rect 3712 10198 3740 10696
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 3068 8922 3096 9930
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9722 3648 9862
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3422 9616 3478 9625
rect 3422 9551 3424 9560
rect 3476 9551 3478 9560
rect 3424 9522 3476 9528
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3169 9276 3477 9285
rect 3169 9274 3175 9276
rect 3231 9274 3255 9276
rect 3311 9274 3335 9276
rect 3391 9274 3415 9276
rect 3471 9274 3477 9276
rect 3231 9222 3233 9274
rect 3413 9222 3415 9274
rect 3169 9220 3175 9222
rect 3231 9220 3255 9222
rect 3311 9220 3335 9222
rect 3391 9220 3415 9222
rect 3471 9220 3477 9222
rect 3169 9211 3477 9220
rect 3240 8968 3292 8974
rect 3068 8894 3188 8922
rect 3240 8910 3292 8916
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 6798 3004 8230
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6361 3004 6598
rect 2962 6352 3018 6361
rect 2962 6287 3018 6296
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 5914 2912 6122
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2976 5778 3004 6054
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5234 2912 5510
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2884 4758 2912 5170
rect 2976 4826 3004 5170
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2962 4176 3018 4185
rect 2780 4140 2832 4146
rect 2962 4111 3018 4120
rect 2780 4082 2832 4088
rect 2976 3738 3004 4111
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2976 3602 3004 3674
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 3068 3534 3096 8774
rect 3160 8566 3188 8894
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3252 8294 3280 8910
rect 3528 8634 3556 9318
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3169 8188 3477 8197
rect 3169 8186 3175 8188
rect 3231 8186 3255 8188
rect 3311 8186 3335 8188
rect 3391 8186 3415 8188
rect 3471 8186 3477 8188
rect 3231 8134 3233 8186
rect 3413 8134 3415 8186
rect 3169 8132 3175 8134
rect 3231 8132 3255 8134
rect 3311 8132 3335 8134
rect 3391 8132 3415 8134
rect 3471 8132 3477 8134
rect 3169 8123 3477 8132
rect 3422 7984 3478 7993
rect 3422 7919 3478 7928
rect 3436 7478 3464 7919
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3528 7206 3556 8570
rect 3620 8566 3648 9046
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3620 7886 3648 8502
rect 3712 8498 3740 10134
rect 3804 9926 3832 10764
rect 4172 10674 4200 11154
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3988 9926 4016 10542
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4080 10441 4108 10474
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3829 9820 4137 9829
rect 3829 9818 3835 9820
rect 3891 9818 3915 9820
rect 3971 9818 3995 9820
rect 4051 9818 4075 9820
rect 4131 9818 4137 9820
rect 3891 9766 3893 9818
rect 4073 9766 4075 9818
rect 3829 9764 3835 9766
rect 3891 9764 3915 9766
rect 3971 9764 3995 9766
rect 4051 9764 4075 9766
rect 4131 9764 4137 9766
rect 3829 9755 4137 9764
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3804 9178 3832 9658
rect 4172 9625 4200 9998
rect 4158 9616 4214 9625
rect 4068 9580 4120 9586
rect 4158 9551 4214 9560
rect 4068 9522 4120 9528
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 4080 8820 4108 9522
rect 4264 9217 4292 12174
rect 4356 12102 4384 13790
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4250 9208 4306 9217
rect 4160 9172 4212 9178
rect 4356 9178 4384 12038
rect 4448 11801 4476 13466
rect 4540 13394 4568 14962
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4632 14618 4660 14758
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4434 11792 4490 11801
rect 4434 11727 4490 11736
rect 4250 9143 4306 9152
rect 4344 9172 4396 9178
rect 4160 9114 4212 9120
rect 4344 9114 4396 9120
rect 4172 9024 4200 9114
rect 4172 8996 4384 9024
rect 4250 8936 4306 8945
rect 4250 8871 4306 8880
rect 4080 8792 4200 8820
rect 3829 8732 4137 8741
rect 3829 8730 3835 8732
rect 3891 8730 3915 8732
rect 3971 8730 3995 8732
rect 4051 8730 4075 8732
rect 4131 8730 4137 8732
rect 3891 8678 3893 8730
rect 4073 8678 4075 8730
rect 3829 8676 3835 8678
rect 3891 8676 3915 8678
rect 3971 8676 3995 8678
rect 4051 8676 4075 8678
rect 4131 8676 4137 8678
rect 3829 8667 4137 8676
rect 4172 8616 4200 8792
rect 4080 8588 4200 8616
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3712 7546 3740 8230
rect 4080 7834 4108 8588
rect 4080 7806 4200 7834
rect 3829 7644 4137 7653
rect 3829 7642 3835 7644
rect 3891 7642 3915 7644
rect 3971 7642 3995 7644
rect 4051 7642 4075 7644
rect 4131 7642 4137 7644
rect 3891 7590 3893 7642
rect 4073 7590 4075 7642
rect 3829 7588 3835 7590
rect 3891 7588 3915 7590
rect 3971 7588 3995 7590
rect 4051 7588 4075 7590
rect 4131 7588 4137 7590
rect 3829 7579 4137 7588
rect 3700 7540 3752 7546
rect 4172 7528 4200 7806
rect 3700 7482 3752 7488
rect 4080 7500 4200 7528
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6225 3464 6598
rect 3422 6216 3478 6225
rect 3422 6151 3478 6160
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 3528 5030 3556 7142
rect 4080 6882 4108 7500
rect 4080 6854 4200 6882
rect 4066 6760 4122 6769
rect 3608 6724 3660 6730
rect 4066 6695 4068 6704
rect 3608 6666 3660 6672
rect 4120 6695 4122 6704
rect 4068 6666 4120 6672
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3344 4282 3372 4490
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3528 3942 3556 4966
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3620 3194 3648 6666
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3712 6186 3740 6598
rect 3829 6556 4137 6565
rect 3829 6554 3835 6556
rect 3891 6554 3915 6556
rect 3971 6554 3995 6556
rect 4051 6554 4075 6556
rect 4131 6554 4137 6556
rect 3891 6502 3893 6554
rect 4073 6502 4075 6554
rect 3829 6500 3835 6502
rect 3891 6500 3915 6502
rect 3971 6500 3995 6502
rect 4051 6500 4075 6502
rect 4131 6500 4137 6502
rect 3829 6491 4137 6500
rect 4172 6440 4200 6854
rect 3804 6412 4200 6440
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3804 5658 3832 6412
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 3712 5630 3832 5658
rect 4172 5642 4200 6258
rect 4264 6254 4292 8871
rect 4356 7886 4384 8996
rect 4448 8974 4476 11727
rect 4540 11150 4568 13330
rect 4632 13138 4660 14554
rect 4710 14240 4766 14249
rect 4710 14175 4766 14184
rect 4724 13258 4752 14175
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4632 13110 4752 13138
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4632 11762 4660 12582
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4618 11656 4674 11665
rect 4724 11626 4752 13110
rect 4618 11591 4674 11600
rect 4712 11620 4764 11626
rect 4632 11354 4660 11591
rect 4712 11562 4764 11568
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4526 10840 4582 10849
rect 4632 10810 4660 11290
rect 4710 11112 4766 11121
rect 4710 11047 4766 11056
rect 4526 10775 4582 10784
rect 4620 10804 4672 10810
rect 4540 10062 4568 10775
rect 4620 10746 4672 10752
rect 4724 10690 4752 11047
rect 4816 10810 4844 15302
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 4896 13864 4948 13870
rect 4894 13832 4896 13841
rect 4948 13832 4950 13841
rect 4894 13767 4950 13776
rect 5000 13716 5028 14962
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 4908 13688 5028 13716
rect 4908 12209 4936 13688
rect 5092 13546 5120 14826
rect 5184 13734 5212 15846
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5000 13518 5120 13546
rect 4894 12200 4950 12209
rect 4894 12135 4950 12144
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4632 10662 4752 10690
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4540 9518 4568 9998
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4540 8838 4568 9318
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4526 8256 4582 8265
rect 4526 8191 4582 8200
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7750 4384 7822
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4342 7032 4398 7041
rect 4342 6967 4398 6976
rect 4356 6798 4384 6967
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4356 6186 4384 6734
rect 4540 6390 4568 8191
rect 4632 7313 4660 10662
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 8129 4752 9862
rect 4710 8120 4766 8129
rect 4710 8055 4766 8064
rect 4618 7304 4674 7313
rect 4618 7239 4674 7248
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4160 5636 4212 5642
rect 3712 3670 3740 5630
rect 4160 5578 4212 5584
rect 3829 5468 4137 5477
rect 3829 5466 3835 5468
rect 3891 5466 3915 5468
rect 3971 5466 3995 5468
rect 4051 5466 4075 5468
rect 4131 5466 4137 5468
rect 3891 5414 3893 5466
rect 4073 5414 4075 5466
rect 3829 5412 3835 5414
rect 3891 5412 3915 5414
rect 3971 5412 3995 5414
rect 4051 5412 4075 5414
rect 4131 5412 4137 5414
rect 3829 5403 4137 5412
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4172 5273 4200 5306
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 4158 5264 4214 5273
rect 4158 5199 4214 5208
rect 3896 4758 3924 5199
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4826 4200 4966
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 4264 4622 4292 5306
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 3829 4380 4137 4389
rect 3829 4378 3835 4380
rect 3891 4378 3915 4380
rect 3971 4378 3995 4380
rect 4051 4378 4075 4380
rect 4131 4378 4137 4380
rect 3891 4326 3893 4378
rect 4073 4326 4075 4378
rect 3829 4324 3835 4326
rect 3891 4324 3915 4326
rect 3971 4324 3995 4326
rect 4051 4324 4075 4326
rect 4131 4324 4137 4326
rect 3829 4315 4137 4324
rect 4356 4282 4384 4558
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4282 4476 4422
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4436 4072 4488 4078
rect 4434 4040 4436 4049
rect 4488 4040 4490 4049
rect 4434 3975 4490 3984
rect 4448 3738 4476 3975
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 4434 3496 4490 3505
rect 4434 3431 4490 3440
rect 4448 3398 4476 3431
rect 4540 3398 4568 6326
rect 4724 5914 4752 8055
rect 4816 7886 4844 10202
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7274 4844 7822
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4908 6186 4936 11494
rect 5000 9994 5028 13518
rect 5080 13184 5132 13190
rect 5078 13152 5080 13161
rect 5132 13152 5134 13161
rect 5078 13087 5134 13096
rect 5184 13002 5212 13670
rect 5276 13569 5304 16458
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5460 15910 5488 16390
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5354 15056 5410 15065
rect 5354 14991 5356 15000
rect 5408 14991 5410 15000
rect 5356 14962 5408 14968
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5262 13560 5318 13569
rect 5262 13495 5318 13504
rect 5092 12974 5212 13002
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 5000 9586 5028 9930
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 5000 8294 5028 9386
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 5000 6066 5028 8230
rect 5092 7886 5120 12974
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5184 12617 5212 12786
rect 5170 12608 5226 12617
rect 5170 12543 5226 12552
rect 5368 12442 5396 14010
rect 5460 13705 5488 15846
rect 5446 13696 5502 13705
rect 5446 13631 5502 13640
rect 5446 13560 5502 13569
rect 5446 13495 5502 13504
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5368 12238 5396 12378
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5172 12096 5224 12102
rect 5460 12073 5488 13495
rect 5552 12306 5580 16594
rect 5644 16250 5672 17070
rect 6012 17066 6040 17138
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5828 16697 5856 16730
rect 5814 16688 5870 16697
rect 5814 16623 5870 16632
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5920 16114 5948 16934
rect 6012 16794 6040 17002
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5828 15502 5856 15846
rect 5816 15496 5868 15502
rect 5920 15473 5948 16050
rect 5998 15600 6054 15609
rect 5998 15535 6054 15544
rect 5816 15438 5868 15444
rect 5906 15464 5962 15473
rect 5906 15399 5962 15408
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5906 15056 5962 15065
rect 5736 14414 5764 15030
rect 5906 14991 5962 15000
rect 5920 14958 5948 14991
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5736 13258 5764 14350
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5172 12038 5224 12044
rect 5446 12064 5502 12073
rect 5184 11393 5212 12038
rect 5446 11999 5502 12008
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5170 11384 5226 11393
rect 5170 11319 5226 11328
rect 5276 11200 5304 11562
rect 5368 11558 5396 11698
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5184 11172 5304 11200
rect 5184 10849 5212 11172
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5170 10840 5226 10849
rect 5276 10810 5304 11018
rect 5170 10775 5226 10784
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5080 7880 5132 7886
rect 5184 7857 5212 10542
rect 5080 7822 5132 7828
rect 5170 7848 5226 7857
rect 5170 7783 5226 7792
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5092 6905 5120 7346
rect 5078 6896 5134 6905
rect 5078 6831 5134 6840
rect 5170 6760 5226 6769
rect 5170 6695 5226 6704
rect 5184 6458 5212 6695
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5172 6316 5224 6322
rect 4908 6038 5028 6066
rect 5092 6276 5172 6304
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4816 4622 4844 5238
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 3829 3292 4137 3301
rect 3829 3290 3835 3292
rect 3891 3290 3915 3292
rect 3971 3290 3995 3292
rect 4051 3290 4075 3292
rect 4131 3290 4137 3292
rect 3891 3238 3893 3290
rect 4073 3238 4075 3290
rect 3829 3236 3835 3238
rect 3891 3236 3915 3238
rect 3971 3236 3995 3238
rect 4051 3236 4075 3238
rect 4131 3236 4137 3238
rect 3829 3227 4137 3236
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 1872 2746 1992 2774
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 940 2576 992 2582
rect 940 2518 992 2524
rect 1872 2446 1900 2746
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 848 2372 900 2378
rect 848 2314 900 2320
rect 572 1896 624 1902
rect 572 1838 624 1844
rect 860 1601 888 2314
rect 2148 2145 2176 2994
rect 3160 2922 3188 3130
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 4448 2650 4476 3334
rect 4540 3194 4568 3334
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4816 2446 4844 4558
rect 4908 4146 4936 6038
rect 5092 5574 5120 6276
rect 5172 6258 5224 6264
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5000 4826 5028 4966
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4988 4616 5040 4622
rect 4986 4584 4988 4593
rect 5184 4593 5212 5578
rect 5040 4584 5042 4593
rect 4986 4519 5042 4528
rect 5170 4584 5226 4593
rect 5170 4519 5226 4528
rect 5276 4486 5304 10746
rect 5368 5098 5396 11494
rect 5552 10849 5580 11630
rect 5538 10840 5594 10849
rect 5448 10804 5500 10810
rect 5538 10775 5594 10784
rect 5448 10746 5500 10752
rect 5460 10266 5488 10746
rect 5552 10266 5580 10775
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5552 9926 5580 9998
rect 5448 9920 5500 9926
rect 5446 9888 5448 9897
rect 5540 9920 5592 9926
rect 5500 9888 5502 9897
rect 5540 9862 5592 9868
rect 5446 9823 5502 9832
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5460 8974 5488 9114
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3194 4936 4082
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2134 2136 2190 2145
rect 2134 2071 2190 2080
rect 846 1592 902 1601
rect 846 1527 902 1536
rect 2792 785 2820 2314
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 2884 105 2912 2382
rect 5276 2310 5304 4422
rect 5368 3398 5396 5034
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 3194 5396 3334
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5460 3058 5488 7754
rect 5552 5710 5580 9862
rect 5644 9654 5672 13126
rect 5736 12646 5764 13194
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 11082 5764 12582
rect 5816 12164 5868 12170
rect 5816 12106 5868 12112
rect 5828 11354 5856 12106
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5736 10742 5764 11018
rect 5814 10976 5870 10985
rect 5814 10911 5870 10920
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5644 9042 5672 9590
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5644 8566 5672 8842
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5644 7993 5672 8502
rect 5630 7984 5686 7993
rect 5630 7919 5686 7928
rect 5644 6730 5672 7919
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5644 6497 5672 6666
rect 5630 6488 5686 6497
rect 5630 6423 5686 6432
rect 5632 6384 5684 6390
rect 5736 6372 5764 9862
rect 5828 7478 5856 10911
rect 5920 10470 5948 14758
rect 6012 13258 6040 15535
rect 6196 14618 6224 17614
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6564 16998 6592 17138
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6656 16454 6684 16526
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6472 15162 6500 16050
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6276 15020 6328 15026
rect 6328 14980 6408 15008
rect 6276 14962 6328 14968
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6104 13802 6132 13942
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6196 13569 6224 14554
rect 6274 13832 6330 13841
rect 6274 13767 6330 13776
rect 6182 13560 6238 13569
rect 6182 13495 6238 13504
rect 6288 13394 6316 13767
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6104 13002 6132 13194
rect 6104 12974 6224 13002
rect 6196 12850 6224 12974
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6092 12640 6144 12646
rect 6090 12608 6092 12617
rect 6144 12608 6146 12617
rect 6090 12543 6146 12552
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6012 11286 6040 12242
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5920 7936 5948 10202
rect 6012 8634 6040 11086
rect 6104 9330 6132 11494
rect 6196 10062 6224 12786
rect 6288 12102 6316 13330
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6288 10588 6316 11222
rect 6380 10742 6408 14980
rect 6472 14958 6500 15098
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14414 6500 14758
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6472 10810 6500 12786
rect 6564 12186 6592 15030
rect 6656 14260 6684 16390
rect 6748 14890 6776 18119
rect 15382 18048 15438 18057
rect 15382 17983 15438 17992
rect 8022 17776 8078 17785
rect 8022 17711 8078 17720
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 6826 17368 6882 17377
rect 7392 17338 7420 17546
rect 7654 17368 7710 17377
rect 6826 17303 6828 17312
rect 6880 17303 6882 17312
rect 7380 17332 7432 17338
rect 6828 17274 6880 17280
rect 7654 17303 7710 17312
rect 7380 17274 7432 17280
rect 7564 17264 7616 17270
rect 7286 17232 7342 17241
rect 7196 17196 7248 17202
rect 7286 17167 7342 17176
rect 7392 17212 7564 17218
rect 7392 17206 7616 17212
rect 7392 17190 7604 17206
rect 7668 17202 7696 17303
rect 7656 17196 7708 17202
rect 7196 17138 7248 17144
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6840 15881 6868 15982
rect 6932 15978 6960 16730
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6826 15872 6882 15881
rect 6826 15807 6882 15816
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6840 15162 6868 15506
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6840 14346 6868 15098
rect 6932 15026 6960 15642
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 7116 14618 7144 16934
rect 7208 16289 7236 17138
rect 7300 16794 7328 17167
rect 7392 16998 7420 17190
rect 7656 17138 7708 17144
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7608 16892 7916 16901
rect 7608 16890 7614 16892
rect 7670 16890 7694 16892
rect 7750 16890 7774 16892
rect 7830 16890 7854 16892
rect 7910 16890 7916 16892
rect 7670 16838 7672 16890
rect 7852 16838 7854 16890
rect 7608 16836 7614 16838
rect 7670 16836 7694 16838
rect 7750 16836 7774 16838
rect 7830 16836 7854 16838
rect 7910 16836 7916 16838
rect 7608 16827 7916 16836
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7286 16552 7342 16561
rect 7286 16487 7342 16496
rect 7194 16280 7250 16289
rect 7194 16215 7250 16224
rect 7300 15570 7328 16487
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7392 15570 7420 15846
rect 7608 15804 7916 15813
rect 7608 15802 7614 15804
rect 7670 15802 7694 15804
rect 7750 15802 7774 15804
rect 7830 15802 7854 15804
rect 7910 15802 7916 15804
rect 7670 15750 7672 15802
rect 7852 15750 7854 15802
rect 7608 15748 7614 15750
rect 7670 15748 7694 15750
rect 7750 15748 7774 15750
rect 7830 15748 7854 15750
rect 7910 15748 7916 15750
rect 7608 15739 7916 15748
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7300 15094 7328 15506
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7288 14952 7340 14958
rect 7392 14940 7420 15506
rect 7340 14912 7420 14940
rect 7472 14952 7524 14958
rect 7288 14894 7340 14900
rect 7944 14929 7972 15846
rect 8036 15162 8064 17711
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 14370 17640 14426 17649
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 8268 17436 8576 17445
rect 8268 17434 8274 17436
rect 8330 17434 8354 17436
rect 8410 17434 8434 17436
rect 8490 17434 8514 17436
rect 8570 17434 8576 17436
rect 8330 17382 8332 17434
rect 8512 17382 8514 17434
rect 8268 17380 8274 17382
rect 8330 17380 8354 17382
rect 8410 17380 8434 17382
rect 8490 17380 8514 17382
rect 8570 17380 8576 17382
rect 8268 17371 8576 17380
rect 12707 17436 13015 17445
rect 12707 17434 12713 17436
rect 12769 17434 12793 17436
rect 12849 17434 12873 17436
rect 12929 17434 12953 17436
rect 13009 17434 13015 17436
rect 12769 17382 12771 17434
rect 12951 17382 12953 17434
rect 12707 17380 12713 17382
rect 12769 17380 12793 17382
rect 12849 17380 12873 17382
rect 12929 17380 12953 17382
rect 13009 17380 13015 17382
rect 12707 17371 13015 17380
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8404 16998 8432 17070
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16697 8432 16934
rect 8390 16688 8446 16697
rect 8390 16623 8446 16632
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16522 8524 16594
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8268 16348 8576 16357
rect 8268 16346 8274 16348
rect 8330 16346 8354 16348
rect 8410 16346 8434 16348
rect 8490 16346 8514 16348
rect 8570 16346 8576 16348
rect 8330 16294 8332 16346
rect 8512 16294 8514 16346
rect 8268 16292 8274 16294
rect 8330 16292 8354 16294
rect 8410 16292 8434 16294
rect 8490 16292 8514 16294
rect 8570 16292 8576 16294
rect 8268 16283 8576 16292
rect 8680 16114 8708 16526
rect 8772 16114 8800 17070
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8864 16114 8892 16934
rect 9140 16658 9168 16934
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8482 16008 8538 16017
rect 8772 15978 8800 16050
rect 8482 15943 8484 15952
rect 8536 15943 8538 15952
rect 8760 15972 8812 15978
rect 8484 15914 8536 15920
rect 8760 15914 8812 15920
rect 8208 15904 8260 15910
rect 8206 15872 8208 15881
rect 8260 15872 8262 15881
rect 8206 15807 8262 15816
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15366 8340 15506
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8268 15260 8576 15269
rect 8268 15258 8274 15260
rect 8330 15258 8354 15260
rect 8410 15258 8434 15260
rect 8490 15258 8514 15260
rect 8570 15258 8576 15260
rect 8330 15206 8332 15258
rect 8512 15206 8514 15258
rect 8268 15204 8274 15206
rect 8330 15204 8354 15206
rect 8410 15204 8434 15206
rect 8490 15204 8514 15206
rect 8570 15204 8576 15206
rect 8268 15195 8576 15204
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8392 15156 8444 15162
rect 8680 15144 8708 15302
rect 8444 15116 8708 15144
rect 8392 15098 8444 15104
rect 8128 15042 8156 15098
rect 8772 15076 8800 15914
rect 8864 15881 8892 16050
rect 8850 15872 8906 15881
rect 8850 15807 8906 15816
rect 8680 15048 8800 15076
rect 8036 15026 8156 15042
rect 8312 15026 8616 15042
rect 8024 15020 8156 15026
rect 8076 15014 8156 15020
rect 8300 15020 8628 15026
rect 8024 14962 8076 14968
rect 8352 15014 8576 15020
rect 8300 14962 8352 14968
rect 8576 14962 8628 14968
rect 7472 14894 7524 14900
rect 7930 14920 7986 14929
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6736 14272 6788 14278
rect 6656 14232 6736 14260
rect 6736 14214 6788 14220
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6748 13326 6776 14214
rect 6932 14006 6960 14214
rect 7116 14113 7144 14554
rect 7102 14104 7158 14113
rect 7102 14039 7158 14048
rect 7116 14006 7144 14039
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6918 13696 6974 13705
rect 6918 13631 6974 13640
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 13190 6776 13262
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6644 12640 6696 12646
rect 6932 12594 6960 13631
rect 6644 12582 6696 12588
rect 6656 12374 6684 12582
rect 6840 12566 6960 12594
rect 6840 12434 6868 12566
rect 7024 12458 7052 13806
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 6748 12406 6868 12434
rect 6932 12430 7052 12458
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6564 12158 6684 12186
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11218 6592 12038
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 6288 10560 6408 10588
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6196 9489 6224 9522
rect 6182 9480 6238 9489
rect 6182 9415 6238 9424
rect 6104 9302 6224 9330
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6104 8362 6132 9114
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6196 8090 6224 9302
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 5920 7908 6132 7936
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5684 6344 5764 6372
rect 5632 6326 5684 6332
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5538 5536 5594 5545
rect 5538 5471 5594 5480
rect 5552 4214 5580 5471
rect 5736 5234 5764 6344
rect 5828 6254 5856 7414
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5920 5574 5948 7686
rect 6012 6186 6040 7754
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6012 5710 6040 5850
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 6104 5273 6132 7908
rect 6288 6984 6316 10066
rect 6380 8090 6408 10560
rect 6458 10432 6514 10441
rect 6458 10367 6514 10376
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6288 6956 6408 6984
rect 6274 6896 6330 6905
rect 6274 6831 6330 6840
rect 6288 5914 6316 6831
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6380 5778 6408 6956
rect 6472 5914 6500 10367
rect 6564 10130 6592 10950
rect 6656 10810 6684 12158
rect 6748 10985 6776 12406
rect 6826 12064 6882 12073
rect 6826 11999 6882 12008
rect 6840 11762 6868 11999
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6840 11558 6868 11698
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6734 10976 6790 10985
rect 6734 10911 6790 10920
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6642 10704 6698 10713
rect 6642 10639 6698 10648
rect 6736 10668 6788 10674
rect 6656 10266 6684 10639
rect 6736 10610 6788 10616
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6642 10160 6698 10169
rect 6552 10124 6604 10130
rect 6642 10095 6698 10104
rect 6552 10066 6604 10072
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6564 6458 6592 9590
rect 6656 9518 6684 10095
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 6458 6684 9318
rect 6748 6866 6776 10610
rect 6840 7750 6868 11290
rect 6932 10033 6960 12430
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6918 9480 6974 9489
rect 6918 9415 6974 9424
rect 6932 9178 6960 9415
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7024 9110 7052 12174
rect 7116 11898 7144 13738
rect 7300 13682 7328 14894
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7208 13654 7328 13682
rect 7208 12170 7236 13654
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7300 11694 7328 12310
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7300 11354 7328 11630
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7286 11112 7342 11121
rect 7286 11047 7288 11056
rect 7340 11047 7342 11056
rect 7288 11018 7340 11024
rect 7392 10742 7420 14486
rect 7484 13938 7512 14894
rect 7930 14855 7986 14864
rect 7608 14716 7916 14725
rect 7608 14714 7614 14716
rect 7670 14714 7694 14716
rect 7750 14714 7774 14716
rect 7830 14714 7854 14716
rect 7910 14714 7916 14716
rect 7670 14662 7672 14714
rect 7852 14662 7854 14714
rect 7608 14660 7614 14662
rect 7670 14660 7694 14662
rect 7750 14660 7774 14662
rect 7830 14660 7854 14662
rect 7910 14660 7916 14662
rect 7608 14651 7916 14660
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7472 13728 7524 13734
rect 7576 13716 7604 14350
rect 8036 14074 8064 14962
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8128 14521 8156 14894
rect 8220 14657 8248 14894
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8206 14648 8262 14657
rect 8206 14583 8262 14592
rect 8496 14521 8524 14758
rect 8114 14512 8170 14521
rect 8114 14447 8170 14456
rect 8482 14512 8538 14521
rect 8482 14447 8538 14456
rect 8116 14408 8168 14414
rect 8680 14396 8708 15048
rect 8956 15026 8984 16594
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 16289 9168 16390
rect 9126 16280 9182 16289
rect 9232 16266 9260 17274
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 12164 17264 12216 17270
rect 12532 17264 12584 17270
rect 12164 17206 12216 17212
rect 12346 17232 12402 17241
rect 9416 16969 9444 17206
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 9402 16960 9458 16969
rect 9402 16895 9458 16904
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9312 16584 9364 16590
rect 9508 16572 9536 16662
rect 9364 16544 9536 16572
rect 9312 16526 9364 16532
rect 9232 16238 9352 16266
rect 9126 16215 9182 16224
rect 9220 16176 9272 16182
rect 9220 16118 9272 16124
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 8852 15020 8904 15026
rect 8772 14980 8852 15008
rect 8772 14550 8800 14980
rect 8852 14962 8904 14968
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8956 14550 8984 14962
rect 9048 14929 9076 16050
rect 9140 16017 9168 16050
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 9126 15328 9182 15337
rect 9126 15263 9182 15272
rect 9034 14920 9090 14929
rect 9034 14855 9090 14864
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 8944 14408 8996 14414
rect 8680 14368 8800 14396
rect 8116 14350 8168 14356
rect 8128 14249 8156 14350
rect 8114 14240 8170 14249
rect 8772 14226 8800 14368
rect 8944 14350 8996 14356
rect 8772 14198 8892 14226
rect 8114 14175 8170 14184
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 7524 13688 7604 13716
rect 8022 13696 8078 13705
rect 7472 13670 7524 13676
rect 7484 13462 7512 13670
rect 7608 13628 7916 13637
rect 8022 13631 8078 13640
rect 7608 13626 7614 13628
rect 7670 13626 7694 13628
rect 7750 13626 7774 13628
rect 7830 13626 7854 13628
rect 7910 13626 7916 13628
rect 7670 13574 7672 13626
rect 7852 13574 7854 13626
rect 7608 13572 7614 13574
rect 7670 13572 7694 13574
rect 7750 13572 7774 13574
rect 7830 13572 7854 13574
rect 7910 13572 7916 13574
rect 7608 13563 7916 13572
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 7484 12782 7512 13398
rect 8036 13394 8064 13631
rect 8128 13462 8156 14175
rect 8268 14172 8576 14181
rect 8268 14170 8274 14172
rect 8330 14170 8354 14172
rect 8410 14170 8434 14172
rect 8490 14170 8514 14172
rect 8570 14170 8576 14172
rect 8330 14118 8332 14170
rect 8512 14118 8514 14170
rect 8268 14116 8274 14118
rect 8330 14116 8354 14118
rect 8410 14116 8434 14118
rect 8490 14116 8514 14118
rect 8570 14116 8576 14118
rect 8268 14107 8576 14116
rect 8758 13968 8814 13977
rect 8758 13903 8814 13912
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 7562 13016 7618 13025
rect 7562 12951 7618 12960
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7576 12628 7604 12951
rect 7668 12918 7696 13330
rect 8268 13084 8576 13093
rect 8268 13082 8274 13084
rect 8330 13082 8354 13084
rect 8410 13082 8434 13084
rect 8490 13082 8514 13084
rect 8570 13082 8576 13084
rect 8330 13030 8332 13082
rect 8512 13030 8514 13082
rect 8268 13028 8274 13030
rect 8330 13028 8354 13030
rect 8410 13028 8434 13030
rect 8490 13028 8514 13030
rect 8570 13028 8576 13030
rect 8268 13019 8576 13028
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 7484 12600 7604 12628
rect 7932 12640 7984 12646
rect 7484 12424 7512 12600
rect 7932 12582 7984 12588
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7608 12540 7916 12549
rect 7608 12538 7614 12540
rect 7670 12538 7694 12540
rect 7750 12538 7774 12540
rect 7830 12538 7854 12540
rect 7910 12538 7916 12540
rect 7670 12486 7672 12538
rect 7852 12486 7854 12538
rect 7608 12484 7614 12486
rect 7670 12484 7694 12486
rect 7750 12484 7774 12486
rect 7830 12484 7854 12486
rect 7910 12484 7916 12486
rect 7608 12475 7916 12484
rect 7748 12436 7800 12442
rect 7484 12396 7604 12424
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7484 10962 7512 12106
rect 7576 11676 7604 12396
rect 7944 12434 7972 12582
rect 7800 12406 7972 12434
rect 7748 12378 7800 12384
rect 7760 12306 7788 12378
rect 8036 12356 8064 12582
rect 8312 12442 8340 12786
rect 8482 12744 8538 12753
rect 8482 12679 8538 12688
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 7852 12328 8064 12356
rect 8114 12336 8170 12345
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7760 11937 7788 12106
rect 7746 11928 7802 11937
rect 7746 11863 7802 11872
rect 7656 11688 7708 11694
rect 7576 11648 7656 11676
rect 7656 11630 7708 11636
rect 7852 11540 7880 12328
rect 7944 12280 8114 12288
rect 7944 12271 8170 12280
rect 7944 12260 8156 12271
rect 7944 11898 7972 12260
rect 8496 12170 8524 12679
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8022 12064 8078 12073
rect 8022 11999 8078 12008
rect 8036 11898 8064 11999
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7852 11512 8064 11540
rect 7608 11452 7916 11461
rect 7608 11450 7614 11452
rect 7670 11450 7694 11452
rect 7750 11450 7774 11452
rect 7830 11450 7854 11452
rect 7910 11450 7916 11452
rect 7670 11398 7672 11450
rect 7852 11398 7854 11450
rect 7608 11396 7614 11398
rect 7670 11396 7694 11398
rect 7750 11396 7774 11398
rect 7830 11396 7854 11398
rect 7910 11396 7916 11398
rect 7608 11387 7916 11396
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7576 11082 7604 11290
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7668 10985 7696 11086
rect 7654 10976 7710 10985
rect 7484 10934 7597 10962
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7116 10606 7144 10678
rect 7104 10600 7156 10606
rect 7484 10554 7512 10746
rect 7569 10724 7597 10934
rect 7654 10911 7710 10920
rect 7746 10840 7802 10849
rect 7746 10775 7748 10784
rect 7800 10775 7802 10784
rect 7748 10746 7800 10752
rect 7852 10742 7880 11086
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7656 10736 7708 10742
rect 7569 10696 7604 10724
rect 7104 10542 7156 10548
rect 7300 10526 7512 10554
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 9722 7144 10406
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7208 9897 7236 10134
rect 7300 10130 7328 10526
rect 7576 10452 7604 10696
rect 7656 10678 7708 10684
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7668 10470 7696 10678
rect 7484 10424 7604 10452
rect 7656 10464 7708 10470
rect 7378 10296 7434 10305
rect 7378 10231 7434 10240
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7392 10062 7420 10231
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7484 9908 7512 10424
rect 7656 10406 7708 10412
rect 7608 10364 7916 10373
rect 7608 10362 7614 10364
rect 7670 10362 7694 10364
rect 7750 10362 7774 10364
rect 7830 10362 7854 10364
rect 7910 10362 7916 10364
rect 7670 10310 7672 10362
rect 7852 10310 7854 10362
rect 7608 10308 7614 10310
rect 7670 10308 7694 10310
rect 7750 10308 7774 10310
rect 7830 10308 7854 10310
rect 7910 10308 7916 10310
rect 7608 10299 7916 10308
rect 7748 10260 7800 10266
rect 7194 9888 7250 9897
rect 7194 9823 7250 9832
rect 7392 9880 7512 9908
rect 7576 10220 7748 10248
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7208 9602 7236 9823
rect 7116 9586 7236 9602
rect 7104 9580 7236 9586
rect 7156 9574 7236 9580
rect 7104 9522 7156 9528
rect 7196 9512 7248 9518
rect 7392 9500 7420 9880
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7196 9454 7248 9460
rect 7300 9472 7420 9500
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6932 8537 6960 8978
rect 7116 8974 7144 9318
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7208 8906 7236 9454
rect 7300 9024 7328 9472
rect 7484 9432 7512 9658
rect 7576 9654 7604 10220
rect 7748 10202 7800 10208
rect 7654 10024 7710 10033
rect 7654 9959 7710 9968
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7392 9404 7512 9432
rect 7392 9092 7420 9404
rect 7668 9364 7696 9959
rect 7484 9336 7696 9364
rect 7484 9160 7512 9336
rect 7608 9276 7916 9285
rect 7608 9274 7614 9276
rect 7670 9274 7694 9276
rect 7750 9274 7774 9276
rect 7830 9274 7854 9276
rect 7910 9274 7916 9276
rect 7670 9222 7672 9274
rect 7852 9222 7854 9274
rect 7608 9220 7614 9222
rect 7670 9220 7694 9222
rect 7750 9220 7774 9222
rect 7830 9220 7854 9222
rect 7910 9220 7916 9222
rect 7608 9211 7916 9220
rect 7748 9172 7800 9178
rect 7484 9132 7604 9160
rect 7392 9064 7512 9092
rect 7300 8996 7420 9024
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7012 8560 7064 8566
rect 6918 8528 6974 8537
rect 7012 8502 7064 8508
rect 6918 8463 6974 8472
rect 6918 8392 6974 8401
rect 6918 8327 6974 8336
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6932 7002 6960 8327
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 6458 6776 6802
rect 7024 6633 7052 8502
rect 7208 8498 7236 8842
rect 7286 8664 7342 8673
rect 7286 8599 7342 8608
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7102 8120 7158 8129
rect 7102 8055 7104 8064
rect 7156 8055 7158 8064
rect 7104 8026 7156 8032
rect 7102 7984 7158 7993
rect 7102 7919 7158 7928
rect 7010 6624 7066 6633
rect 7010 6559 7066 6568
rect 7010 6488 7066 6497
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6736 6452 6788 6458
rect 7116 6458 7144 7919
rect 7208 6730 7236 8434
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7010 6423 7066 6432
rect 7104 6452 7156 6458
rect 6736 6394 6788 6400
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6656 6202 6684 6394
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6274 5672 6330 5681
rect 6274 5607 6330 5616
rect 6090 5264 6146 5273
rect 5724 5228 5776 5234
rect 6090 5199 6146 5208
rect 5724 5170 5776 5176
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5736 3534 5764 3674
rect 6104 3618 6132 5199
rect 6288 4146 6316 5607
rect 6380 5030 6408 5714
rect 6472 5642 6500 5850
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6564 5114 6592 6190
rect 6656 6174 6868 6202
rect 6840 6118 6868 6174
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6828 6112 6880 6118
rect 6932 6089 6960 6122
rect 6828 6054 6880 6060
rect 6918 6080 6974 6089
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5234 6776 5510
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6472 5086 6592 5114
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6472 4758 6500 5086
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6012 3590 6132 3618
rect 5540 3528 5592 3534
rect 5632 3528 5684 3534
rect 5540 3470 5592 3476
rect 5630 3496 5632 3505
rect 5724 3528 5776 3534
rect 5684 3496 5686 3505
rect 5552 3194 5580 3470
rect 5724 3470 5776 3476
rect 5630 3431 5686 3440
rect 6012 3194 6040 3590
rect 6090 3496 6146 3505
rect 6090 3431 6092 3440
rect 6144 3431 6146 3440
rect 6092 3402 6144 3408
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 6196 2514 6224 3946
rect 6458 3768 6514 3777
rect 6458 3703 6460 3712
rect 6512 3703 6514 3712
rect 6460 3674 6512 3680
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 6288 2990 6316 3402
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6564 2650 6592 4966
rect 6656 4758 6684 5102
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6840 2854 6868 6054
rect 6918 6015 6974 6024
rect 7024 5302 7052 6423
rect 7104 6394 7156 6400
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 7300 4690 7328 8599
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7392 2990 7420 8996
rect 7484 6905 7512 9064
rect 7576 8566 7604 9132
rect 7748 9114 7800 9120
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7760 8401 7788 9114
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 8809 7880 8978
rect 7838 8800 7894 8809
rect 7838 8735 7894 8744
rect 7746 8392 7802 8401
rect 7746 8327 7802 8336
rect 7608 8188 7916 8197
rect 7608 8186 7614 8188
rect 7670 8186 7694 8188
rect 7750 8186 7774 8188
rect 7830 8186 7854 8188
rect 7910 8186 7916 8188
rect 7670 8134 7672 8186
rect 7852 8134 7854 8186
rect 7608 8132 7614 8134
rect 7670 8132 7694 8134
rect 7750 8132 7774 8134
rect 7830 8132 7854 8134
rect 7910 8132 7916 8134
rect 7608 8123 7916 8132
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 7470 6896 7526 6905
rect 7470 6831 7526 6840
rect 7654 6624 7710 6633
rect 7654 6559 7710 6568
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 5574 7512 6190
rect 7668 6186 7696 6559
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7470 5264 7526 5273
rect 7470 5199 7526 5208
rect 7484 4808 7512 5199
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 7484 4780 7604 4808
rect 7576 4622 7604 4780
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 3194 7512 4082
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 7838 3632 7894 3641
rect 7838 3567 7894 3576
rect 7852 3398 7880 3567
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 7484 2650 7512 3130
rect 7944 3126 7972 10950
rect 8036 6066 8064 11512
rect 8128 11150 8156 12106
rect 8268 11996 8576 12005
rect 8268 11994 8274 11996
rect 8330 11994 8354 11996
rect 8410 11994 8434 11996
rect 8490 11994 8514 11996
rect 8570 11994 8576 11996
rect 8330 11942 8332 11994
rect 8512 11942 8514 11994
rect 8268 11940 8274 11942
rect 8330 11940 8354 11942
rect 8410 11940 8434 11942
rect 8490 11940 8514 11942
rect 8570 11940 8576 11942
rect 8268 11931 8576 11940
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8404 11393 8432 11630
rect 8588 11558 8616 11630
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8390 11384 8446 11393
rect 8390 11319 8446 11328
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10470 8156 10950
rect 8268 10908 8576 10917
rect 8268 10906 8274 10908
rect 8330 10906 8354 10908
rect 8410 10906 8434 10908
rect 8490 10906 8514 10908
rect 8570 10906 8576 10908
rect 8330 10854 8332 10906
rect 8512 10854 8514 10906
rect 8268 10852 8274 10854
rect 8330 10852 8354 10854
rect 8410 10852 8434 10854
rect 8490 10852 8514 10854
rect 8570 10852 8576 10854
rect 8268 10843 8576 10852
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8574 10704 8630 10713
rect 8220 10470 8248 10678
rect 8574 10639 8576 10648
rect 8628 10639 8630 10648
rect 8576 10610 8628 10616
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8208 10464 8260 10470
rect 8496 10441 8524 10474
rect 8208 10406 8260 10412
rect 8482 10432 8538 10441
rect 8220 10266 8248 10406
rect 8482 10367 8538 10376
rect 8588 10266 8616 10610
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8298 10160 8354 10169
rect 8128 10118 8298 10146
rect 8128 8673 8156 10118
rect 8298 10095 8354 10104
rect 8208 10056 8260 10062
rect 8206 10024 8208 10033
rect 8260 10024 8262 10033
rect 8206 9959 8262 9968
rect 8268 9820 8576 9829
rect 8268 9818 8274 9820
rect 8330 9818 8354 9820
rect 8410 9818 8434 9820
rect 8490 9818 8514 9820
rect 8570 9818 8576 9820
rect 8330 9766 8332 9818
rect 8512 9766 8514 9818
rect 8268 9764 8274 9766
rect 8330 9764 8354 9766
rect 8410 9764 8434 9766
rect 8490 9764 8514 9766
rect 8570 9764 8576 9766
rect 8268 9755 8576 9764
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8220 9382 8248 9590
rect 8680 9518 8708 13806
rect 8772 13025 8800 13903
rect 8758 13016 8814 13025
rect 8758 12951 8814 12960
rect 8864 12918 8892 14198
rect 8956 13841 8984 14350
rect 9140 13954 9168 15263
rect 9232 15162 9260 16118
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9232 14822 9260 14962
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9048 13926 9168 13954
rect 8942 13832 8998 13841
rect 8942 13767 8998 13776
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 8906 8248 9318
rect 8390 9208 8446 9217
rect 8390 9143 8446 9152
rect 8404 9042 8432 9143
rect 8772 9058 8800 12038
rect 8864 11830 8892 12650
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8864 9897 8892 10134
rect 8850 9888 8906 9897
rect 8850 9823 8906 9832
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8680 9030 8800 9058
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8268 8732 8576 8741
rect 8268 8730 8274 8732
rect 8330 8730 8354 8732
rect 8410 8730 8434 8732
rect 8490 8730 8514 8732
rect 8570 8730 8576 8732
rect 8330 8678 8332 8730
rect 8512 8678 8514 8730
rect 8268 8676 8274 8678
rect 8330 8676 8354 8678
rect 8410 8676 8434 8678
rect 8490 8676 8514 8678
rect 8570 8676 8576 8678
rect 8114 8664 8170 8673
rect 8268 8667 8576 8676
rect 8114 8599 8170 8608
rect 8392 8628 8444 8634
rect 8128 8566 8156 8599
rect 8392 8570 8444 8576
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8114 8392 8170 8401
rect 8114 8327 8170 8336
rect 8128 6390 8156 8327
rect 8404 7886 8432 8570
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8496 8362 8524 8502
rect 8680 8430 8708 9030
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 8498 8800 8910
rect 8864 8566 8892 9454
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8496 7834 8524 8298
rect 8588 8090 8616 8298
rect 8576 8084 8628 8090
rect 8628 8044 8800 8072
rect 8576 8026 8628 8032
rect 8496 7806 8708 7834
rect 8268 7644 8576 7653
rect 8268 7642 8274 7644
rect 8330 7642 8354 7644
rect 8410 7642 8434 7644
rect 8490 7642 8514 7644
rect 8570 7642 8576 7644
rect 8330 7590 8332 7642
rect 8512 7590 8514 7642
rect 8268 7588 8274 7590
rect 8330 7588 8354 7590
rect 8410 7588 8434 7590
rect 8490 7588 8514 7590
rect 8570 7588 8576 7590
rect 8268 7579 8576 7588
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8312 6934 8340 7210
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8680 6798 8708 7806
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8268 6556 8576 6565
rect 8268 6554 8274 6556
rect 8330 6554 8354 6556
rect 8410 6554 8434 6556
rect 8490 6554 8514 6556
rect 8570 6554 8576 6556
rect 8330 6502 8332 6554
rect 8512 6502 8514 6554
rect 8268 6500 8274 6502
rect 8330 6500 8354 6502
rect 8410 6500 8434 6502
rect 8490 6500 8514 6502
rect 8570 6500 8576 6502
rect 8268 6491 8576 6500
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8116 6180 8168 6186
rect 8168 6140 8248 6168
rect 8116 6122 8168 6128
rect 8036 6038 8156 6066
rect 8022 5944 8078 5953
rect 8022 5879 8078 5888
rect 8036 5642 8064 5879
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8024 5160 8076 5166
rect 8022 5128 8024 5137
rect 8076 5128 8078 5137
rect 8022 5063 8078 5072
rect 8022 4856 8078 4865
rect 8022 4791 8078 4800
rect 8036 4457 8064 4791
rect 8022 4448 8078 4457
rect 8022 4383 8078 4392
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 8036 3534 8064 3975
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 8128 3058 8156 6038
rect 8220 5681 8248 6140
rect 8404 5914 8432 6394
rect 8772 6254 8800 8044
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8482 5944 8538 5953
rect 8392 5908 8444 5914
rect 8666 5944 8722 5953
rect 8538 5902 8616 5930
rect 8482 5879 8538 5888
rect 8392 5850 8444 5856
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8206 5672 8262 5681
rect 8496 5642 8524 5782
rect 8588 5778 8616 5902
rect 8666 5879 8722 5888
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8206 5607 8262 5616
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8268 5468 8576 5477
rect 8268 5466 8274 5468
rect 8330 5466 8354 5468
rect 8410 5466 8434 5468
rect 8490 5466 8514 5468
rect 8570 5466 8576 5468
rect 8330 5414 8332 5466
rect 8512 5414 8514 5466
rect 8268 5412 8274 5414
rect 8330 5412 8354 5414
rect 8410 5412 8434 5414
rect 8490 5412 8514 5414
rect 8570 5412 8576 5414
rect 8268 5403 8576 5412
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8496 4758 8524 5102
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8268 4380 8576 4389
rect 8268 4378 8274 4380
rect 8330 4378 8354 4380
rect 8410 4378 8434 4380
rect 8490 4378 8514 4380
rect 8570 4378 8576 4380
rect 8330 4326 8332 4378
rect 8512 4326 8514 4378
rect 8268 4324 8274 4326
rect 8330 4324 8354 4326
rect 8410 4324 8434 4326
rect 8490 4324 8514 4326
rect 8570 4324 8576 4326
rect 8268 4315 8576 4324
rect 8680 3534 8708 5879
rect 8864 4282 8892 8366
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8956 4146 8984 12854
rect 9048 11286 9076 13926
rect 9232 13802 9260 14758
rect 9324 14482 9352 16238
rect 9402 15464 9458 15473
rect 9402 15399 9458 15408
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9416 14278 9444 15399
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9312 14000 9364 14006
rect 9508 13977 9536 16544
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9586 16280 9642 16289
rect 9586 16215 9642 16224
rect 9600 15473 9628 16215
rect 9586 15464 9642 15473
rect 9586 15399 9642 15408
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9312 13942 9364 13948
rect 9494 13968 9550 13977
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9324 13734 9352 13942
rect 9404 13932 9456 13938
rect 9494 13903 9550 13912
rect 9404 13874 9456 13880
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9218 13152 9274 13161
rect 9140 12986 9168 13126
rect 9218 13087 9274 13096
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9232 12617 9260 13087
rect 9218 12608 9274 12617
rect 9218 12543 9274 12552
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9034 10704 9090 10713
rect 9034 10639 9090 10648
rect 9048 8362 9076 10639
rect 9140 9625 9168 12174
rect 9218 11928 9274 11937
rect 9218 11863 9220 11872
rect 9272 11863 9274 11872
rect 9220 11834 9272 11840
rect 9324 11778 9352 13670
rect 9416 13308 9444 13874
rect 9416 13280 9536 13308
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12442 9444 13126
rect 9508 12782 9536 13280
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9416 11898 9444 12378
rect 9496 12232 9548 12238
rect 9600 12220 9628 14282
rect 9692 13870 9720 16526
rect 9784 13870 9812 17138
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9968 14006 9996 15302
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 10060 14521 10088 14894
rect 10046 14512 10102 14521
rect 10152 14482 10180 16526
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 15910 10364 16390
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10244 14521 10272 15574
rect 10230 14512 10286 14521
rect 10046 14447 10102 14456
rect 10140 14476 10192 14482
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9692 13682 9720 13806
rect 9692 13654 9812 13682
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9692 12850 9720 13262
rect 9784 13190 9812 13654
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9680 12844 9732 12850
rect 9732 12804 9812 12832
rect 9680 12786 9732 12792
rect 9784 12764 9812 12804
rect 9864 12776 9916 12782
rect 9784 12736 9864 12764
rect 9678 12472 9734 12481
rect 9678 12407 9734 12416
rect 9548 12192 9628 12220
rect 9496 12174 9548 12180
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9220 11756 9272 11762
rect 9324 11750 9444 11778
rect 9220 11698 9272 11704
rect 9232 11558 9260 11698
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9126 9616 9182 9625
rect 9126 9551 9182 9560
rect 9140 8401 9168 9551
rect 9232 8974 9260 11494
rect 9324 11150 9352 11494
rect 9416 11286 9444 11750
rect 9600 11665 9628 12038
rect 9586 11656 9642 11665
rect 9586 11591 9642 11600
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9416 10810 9444 11222
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9402 10704 9458 10713
rect 9402 10639 9458 10648
rect 9310 10296 9366 10305
rect 9310 10231 9312 10240
rect 9364 10231 9366 10240
rect 9312 10202 9364 10208
rect 9324 10062 9352 10202
rect 9416 10198 9444 10639
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9416 9722 9444 10134
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9324 8616 9352 9522
rect 9232 8588 9352 8616
rect 9126 8392 9182 8401
rect 9036 8356 9088 8362
rect 9126 8327 9182 8336
rect 9036 8298 9088 8304
rect 9126 8256 9182 8265
rect 9126 8191 9182 8200
rect 9036 7744 9088 7750
rect 9034 7712 9036 7721
rect 9088 7712 9090 7721
rect 9034 7647 9090 7656
rect 9034 7440 9090 7449
rect 9034 7375 9090 7384
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9048 4010 9076 7375
rect 9140 6390 9168 8191
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9232 5370 9260 8588
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9324 6866 9352 8434
rect 9416 8129 9444 9658
rect 9508 8634 9536 11154
rect 9600 11082 9628 11591
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9588 10804 9640 10810
rect 9692 10792 9720 12407
rect 9784 11150 9812 12736
rect 9864 12718 9916 12724
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9876 12442 9904 12582
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9640 10764 9720 10792
rect 9588 10746 9640 10752
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9600 9926 9628 10610
rect 9692 10266 9720 10610
rect 9770 10296 9826 10305
rect 9680 10260 9732 10266
rect 9770 10231 9826 10240
rect 9680 10202 9732 10208
rect 9692 9994 9720 10202
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9692 9586 9720 9658
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9680 9444 9732 9450
rect 9784 9432 9812 10231
rect 9732 9404 9812 9432
rect 9680 9386 9732 9392
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9081 9628 9318
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9586 9072 9642 9081
rect 9586 9007 9642 9016
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9600 8634 9628 8910
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9402 8120 9458 8129
rect 9402 8055 9458 8064
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9496 7948 9548 7954
rect 9548 7908 9628 7936
rect 9496 7890 9548 7896
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9324 6458 9352 6802
rect 9416 6458 9444 7890
rect 9600 7478 9628 7908
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9600 7342 9628 7414
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9494 6488 9550 6497
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9404 6452 9456 6458
rect 9494 6423 9550 6432
rect 9404 6394 9456 6400
rect 9416 5642 9444 6394
rect 9508 6390 9536 6423
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 4729 9444 5306
rect 9402 4720 9458 4729
rect 9402 4655 9458 4664
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8268 3292 8576 3301
rect 8268 3290 8274 3292
rect 8330 3290 8354 3292
rect 8410 3290 8434 3292
rect 8490 3290 8514 3292
rect 8570 3290 8576 3292
rect 8330 3238 8332 3290
rect 8512 3238 8514 3290
rect 8268 3236 8274 3238
rect 8330 3236 8354 3238
rect 8410 3236 8434 3238
rect 8490 3236 8514 3238
rect 8570 3236 8576 3238
rect 8268 3227 8576 3236
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 3829 2204 4137 2213
rect 3829 2202 3835 2204
rect 3891 2202 3915 2204
rect 3971 2202 3995 2204
rect 4051 2202 4075 2204
rect 4131 2202 4137 2204
rect 3891 2150 3893 2202
rect 4073 2150 4075 2202
rect 3829 2148 3835 2150
rect 3891 2148 3915 2150
rect 3971 2148 3995 2150
rect 4051 2148 4075 2150
rect 4131 2148 4137 2150
rect 3829 2139 4137 2148
rect 7208 1970 7236 2518
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7196 1964 7248 1970
rect 7196 1906 7248 1912
rect 7760 800 7788 2382
rect 8128 2106 8156 2994
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8312 2514 8340 2926
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8680 2446 8708 3334
rect 8772 3058 8800 3606
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2582 8800 2790
rect 8956 2582 8984 2994
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 9048 2446 9076 3334
rect 9600 3058 9628 6598
rect 9692 4690 9720 9114
rect 9784 8974 9812 9404
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9968 8294 9996 13466
rect 10060 12714 10088 14447
rect 10230 14447 10286 14456
rect 10140 14418 10192 14424
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 13258 10180 14214
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10152 13161 10180 13194
rect 10138 13152 10194 13161
rect 10138 13087 10194 13096
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10244 11812 10272 13874
rect 10336 12084 10364 15846
rect 10416 15088 10468 15094
rect 10416 15030 10468 15036
rect 10428 13938 10456 15030
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10428 12986 10456 13466
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10414 12608 10470 12617
rect 10414 12543 10470 12552
rect 10428 12345 10456 12543
rect 10414 12336 10470 12345
rect 10414 12271 10470 12280
rect 10416 12096 10468 12102
rect 10336 12056 10416 12084
rect 10416 12038 10468 12044
rect 10152 11784 10272 11812
rect 10046 11656 10102 11665
rect 10046 11591 10102 11600
rect 10060 10577 10088 11591
rect 10046 10568 10102 10577
rect 10046 10503 10102 10512
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9876 8266 9996 8294
rect 9876 7954 9904 8266
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9772 7744 9824 7750
rect 9956 7744 10008 7750
rect 9824 7704 9904 7732
rect 9772 7686 9824 7692
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9784 7206 9812 7482
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9876 6633 9904 7704
rect 9956 7686 10008 7692
rect 9968 7546 9996 7686
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9862 6624 9918 6633
rect 9862 6559 9918 6568
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9784 5234 9812 6258
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9784 4282 9812 5170
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9692 2446 9720 2926
rect 9876 2922 9904 6559
rect 9968 5794 9996 7210
rect 10060 6390 10088 10406
rect 10152 9217 10180 11784
rect 10322 11520 10378 11529
rect 10322 11455 10378 11464
rect 10336 11200 10364 11455
rect 10428 11268 10456 12038
rect 10520 11393 10548 14758
rect 10506 11384 10562 11393
rect 10506 11319 10562 11328
rect 10428 11240 10548 11268
rect 10336 11172 10456 11200
rect 10230 10704 10286 10713
rect 10230 10639 10286 10648
rect 10244 10606 10272 10639
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 9722 10272 10406
rect 10322 10296 10378 10305
rect 10322 10231 10378 10240
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10230 9616 10286 9625
rect 10230 9551 10286 9560
rect 10244 9518 10272 9551
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10138 9208 10194 9217
rect 10336 9178 10364 10231
rect 10138 9143 10194 9152
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10152 6458 10180 8910
rect 10336 7936 10364 8910
rect 10428 8634 10456 11172
rect 10520 9654 10548 11240
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10520 9518 10548 9590
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10520 9382 10548 9454
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10244 7908 10364 7936
rect 10244 7750 10272 7908
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 9968 5766 10088 5794
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 8268 2204 8576 2213
rect 8268 2202 8274 2204
rect 8330 2202 8354 2204
rect 8410 2202 8434 2204
rect 8490 2202 8514 2204
rect 8570 2202 8576 2204
rect 8330 2150 8332 2202
rect 8512 2150 8514 2202
rect 8268 2148 8274 2150
rect 8330 2148 8354 2150
rect 8410 2148 8434 2150
rect 8490 2148 8514 2150
rect 8570 2148 8576 2150
rect 8268 2139 8576 2148
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 8404 870 8524 898
rect 8404 800 8432 870
rect 2870 96 2926 105
rect 2870 31 2926 40
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 8496 762 8524 870
rect 8680 762 8708 2382
rect 9048 800 9076 2382
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 2038 9260 2246
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9692 800 9720 2382
rect 9968 2310 9996 5646
rect 10060 5273 10088 5766
rect 10046 5264 10102 5273
rect 10046 5199 10102 5208
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10060 3466 10088 3674
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10152 3194 10180 6122
rect 10244 5778 10272 7686
rect 10324 5840 10376 5846
rect 10322 5808 10324 5817
rect 10376 5808 10378 5817
rect 10232 5772 10284 5778
rect 10322 5743 10378 5752
rect 10232 5714 10284 5720
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10152 2922 10180 3130
rect 10140 2916 10192 2922
rect 10140 2858 10192 2864
rect 10244 2650 10272 5170
rect 10322 4176 10378 4185
rect 10322 4111 10378 4120
rect 10336 3194 10364 4111
rect 10428 3738 10456 7754
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 7478 10548 7686
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10520 7002 10548 7414
rect 10612 7410 10640 16186
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10704 9722 10732 14826
rect 10796 14414 10824 16934
rect 10966 16688 11022 16697
rect 10966 16623 11022 16632
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 14249 10824 14350
rect 10782 14240 10838 14249
rect 10782 14175 10838 14184
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10796 10810 10824 13738
rect 10888 13326 10916 15302
rect 10980 15201 11008 16623
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10966 15192 11022 15201
rect 10966 15127 11022 15136
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10980 13326 11008 14554
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10876 12912 10928 12918
rect 11072 12866 11100 16458
rect 11164 12986 11192 17002
rect 11808 16998 11836 17138
rect 12176 17105 12204 17206
rect 12346 17167 12402 17176
rect 12452 17212 12532 17218
rect 12452 17206 12584 17212
rect 12452 17190 12572 17206
rect 12162 17096 12218 17105
rect 12162 17031 12218 17040
rect 12360 17048 12388 17167
rect 12452 17048 12480 17190
rect 12360 17020 12480 17048
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 12047 16892 12355 16901
rect 12047 16890 12053 16892
rect 12109 16890 12133 16892
rect 12189 16890 12213 16892
rect 12269 16890 12293 16892
rect 12349 16890 12355 16892
rect 12109 16838 12111 16890
rect 12291 16838 12293 16890
rect 12047 16836 12053 16838
rect 12109 16836 12133 16838
rect 12189 16836 12213 16838
rect 12269 16836 12293 16838
rect 12349 16836 12355 16838
rect 12047 16827 12355 16836
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11256 16697 11284 16730
rect 11520 16720 11572 16726
rect 11242 16688 11298 16697
rect 11520 16662 11572 16668
rect 11242 16623 11298 16632
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15570 11284 15846
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11256 14618 11284 15370
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11348 14074 11376 15438
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11242 13288 11298 13297
rect 11242 13223 11244 13232
rect 11296 13223 11298 13232
rect 11336 13252 11388 13258
rect 11244 13194 11296 13200
rect 11336 13194 11388 13200
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 10876 12854 10928 12860
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10784 10192 10836 10198
rect 10782 10160 10784 10169
rect 10836 10160 10838 10169
rect 10782 10095 10838 10104
rect 10888 10044 10916 12854
rect 10980 12838 11100 12866
rect 10980 11762 11008 12838
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11060 12232 11112 12238
rect 11058 12200 11060 12209
rect 11112 12200 11114 12209
rect 11058 12135 11114 12144
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11072 11626 11100 12038
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10966 10432 11022 10441
rect 10966 10367 11022 10376
rect 10796 10016 10916 10044
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10704 9042 10732 9114
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 7954 10732 8434
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10704 6780 10732 7890
rect 10796 7290 10824 10016
rect 10980 9994 11008 10367
rect 11072 10198 11100 10950
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 7750 10916 9862
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10980 9110 11008 9658
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 11072 8673 11100 9318
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 11164 8566 11192 12650
rect 11348 12617 11376 13194
rect 11334 12608 11390 12617
rect 11334 12543 11390 12552
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11256 10810 11284 12378
rect 11336 11824 11388 11830
rect 11334 11792 11336 11801
rect 11388 11792 11390 11801
rect 11334 11727 11390 11736
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11354 11376 11494
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11336 10736 11388 10742
rect 11242 10704 11298 10713
rect 11336 10678 11388 10684
rect 11242 10639 11298 10648
rect 11256 9926 11284 10639
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11244 9648 11296 9654
rect 11242 9616 11244 9625
rect 11296 9616 11298 9625
rect 11242 9551 11298 9560
rect 11242 9208 11298 9217
rect 11242 9143 11298 9152
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10796 7262 11008 7290
rect 10784 6792 10836 6798
rect 10704 6752 10784 6780
rect 10784 6734 10836 6740
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10612 5642 10640 6258
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10598 5536 10654 5545
rect 10598 5471 10654 5480
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10336 2446 10364 2926
rect 10612 2650 10640 5471
rect 10704 3534 10732 5714
rect 10796 4214 10824 6734
rect 10980 6225 11008 7262
rect 11072 6662 11100 8298
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7410 11192 7822
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11256 6662 11284 9143
rect 11348 8498 11376 10678
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 8022 11376 8230
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 10966 6216 11022 6225
rect 10966 6151 11022 6160
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 11164 3942 11192 5782
rect 11256 5642 11284 6394
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11348 3738 11376 7686
rect 11440 6458 11468 15030
rect 11532 11354 11560 16662
rect 12084 16590 12112 16730
rect 12256 16720 12308 16726
rect 12452 16708 12480 17020
rect 12308 16680 12480 16708
rect 12256 16662 12308 16668
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11992 16454 12020 16526
rect 13096 16454 13124 17478
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13648 16998 13676 17138
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12530 16280 12586 16289
rect 12530 16215 12532 16224
rect 12584 16215 12586 16224
rect 12532 16186 12584 16192
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11624 15366 11652 15982
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11716 13954 11744 15846
rect 11624 13926 11744 13954
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11532 10606 11560 11290
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11624 10062 11652 13926
rect 11808 13705 11836 16118
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15722 11928 15846
rect 12047 15804 12355 15813
rect 12047 15802 12053 15804
rect 12109 15802 12133 15804
rect 12189 15802 12213 15804
rect 12269 15802 12293 15804
rect 12349 15802 12355 15804
rect 12109 15750 12111 15802
rect 12291 15750 12293 15802
rect 12047 15748 12053 15750
rect 12109 15748 12133 15750
rect 12189 15748 12213 15750
rect 12269 15748 12293 15750
rect 12349 15748 12355 15750
rect 12047 15739 12355 15748
rect 11900 15694 12020 15722
rect 11992 15570 12020 15694
rect 12544 15609 12572 15914
rect 12530 15600 12586 15609
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11980 15564 12032 15570
rect 12530 15535 12586 15544
rect 11980 15506 12032 15512
rect 11900 14958 11928 15506
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12084 15337 12112 15438
rect 12070 15328 12126 15337
rect 12070 15263 12126 15272
rect 12438 15056 12494 15065
rect 12438 14991 12494 15000
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11900 14482 11928 14894
rect 12452 14793 12480 14991
rect 12438 14784 12494 14793
rect 12047 14716 12355 14725
rect 12438 14719 12494 14728
rect 12047 14714 12053 14716
rect 12109 14714 12133 14716
rect 12189 14714 12213 14716
rect 12269 14714 12293 14716
rect 12349 14714 12355 14716
rect 12109 14662 12111 14714
rect 12291 14662 12293 14714
rect 12047 14660 12053 14662
rect 12109 14660 12133 14662
rect 12189 14660 12213 14662
rect 12269 14660 12293 14662
rect 12349 14660 12355 14662
rect 12047 14651 12355 14660
rect 12636 14634 12664 16390
rect 12707 16348 13015 16357
rect 12707 16346 12713 16348
rect 12769 16346 12793 16348
rect 12849 16346 12873 16348
rect 12929 16346 12953 16348
rect 13009 16346 13015 16348
rect 12769 16294 12771 16346
rect 12951 16294 12953 16346
rect 12707 16292 12713 16294
rect 12769 16292 12793 16294
rect 12849 16292 12873 16294
rect 12929 16292 12953 16294
rect 13009 16292 13015 16294
rect 12707 16283 13015 16292
rect 12714 16144 12770 16153
rect 12714 16079 12716 16088
rect 12768 16079 12770 16088
rect 12716 16050 12768 16056
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 13004 15706 13032 15982
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13096 15434 13124 15846
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 12707 15260 13015 15269
rect 12707 15258 12713 15260
rect 12769 15258 12793 15260
rect 12849 15258 12873 15260
rect 12929 15258 12953 15260
rect 13009 15258 13015 15260
rect 12769 15206 12771 15258
rect 12951 15206 12953 15258
rect 12707 15204 12713 15206
rect 12769 15204 12793 15206
rect 12849 15204 12873 15206
rect 12929 15204 12953 15206
rect 13009 15204 13015 15206
rect 12707 15195 13015 15204
rect 12992 15088 13044 15094
rect 13096 15076 13124 15370
rect 13044 15048 13124 15076
rect 12992 15030 13044 15036
rect 12452 14606 12664 14634
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11888 13728 11940 13734
rect 11794 13696 11850 13705
rect 11888 13670 11940 13676
rect 11794 13631 11850 13640
rect 11900 13462 11928 13670
rect 12047 13628 12355 13637
rect 12047 13626 12053 13628
rect 12109 13626 12133 13628
rect 12189 13626 12213 13628
rect 12269 13626 12293 13628
rect 12349 13626 12355 13628
rect 12109 13574 12111 13626
rect 12291 13574 12293 13626
rect 12047 13572 12053 13574
rect 12109 13572 12133 13574
rect 12189 13572 12213 13574
rect 12269 13572 12293 13574
rect 12349 13572 12355 13574
rect 12047 13563 12355 13572
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12268 13326 12296 13398
rect 12072 13320 12124 13326
rect 12070 13288 12072 13297
rect 12256 13320 12308 13326
rect 12124 13288 12126 13297
rect 12256 13262 12308 13268
rect 12070 13223 12126 13232
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11794 12880 11850 12889
rect 11794 12815 11850 12824
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11716 12306 11744 12718
rect 11808 12442 11836 12815
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 11642 11744 12038
rect 11808 11762 11836 12174
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11716 11614 11836 11642
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 10305 11744 10406
rect 11702 10296 11758 10305
rect 11702 10231 11758 10240
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11532 9761 11560 9998
rect 11518 9752 11574 9761
rect 11518 9687 11574 9696
rect 11808 9654 11836 11614
rect 11900 10742 11928 13126
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12176 12782 12204 12922
rect 12164 12776 12216 12782
rect 12268 12753 12296 12922
rect 12164 12718 12216 12724
rect 12254 12744 12310 12753
rect 12254 12679 12310 12688
rect 12047 12540 12355 12549
rect 12047 12538 12053 12540
rect 12109 12538 12133 12540
rect 12189 12538 12213 12540
rect 12269 12538 12293 12540
rect 12349 12538 12355 12540
rect 12109 12486 12111 12538
rect 12291 12486 12293 12538
rect 12047 12484 12053 12486
rect 12109 12484 12133 12486
rect 12189 12484 12213 12486
rect 12269 12484 12293 12486
rect 12349 12484 12355 12486
rect 12047 12475 12355 12484
rect 12452 12434 12480 14606
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12544 13938 12572 14214
rect 12707 14172 13015 14181
rect 12707 14170 12713 14172
rect 12769 14170 12793 14172
rect 12849 14170 12873 14172
rect 12929 14170 12953 14172
rect 13009 14170 13015 14172
rect 12769 14118 12771 14170
rect 12951 14118 12953 14170
rect 12707 14116 12713 14118
rect 12769 14116 12793 14118
rect 12849 14116 12873 14118
rect 12929 14116 12953 14118
rect 13009 14116 13015 14118
rect 12707 14107 13015 14116
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12636 12866 12664 14010
rect 12898 13968 12954 13977
rect 13004 13938 13032 14010
rect 12898 13903 12954 13912
rect 12992 13932 13044 13938
rect 12912 13462 12940 13903
rect 12992 13874 13044 13880
rect 13004 13546 13032 13874
rect 13096 13734 13124 15048
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13004 13518 13124 13546
rect 13280 13530 13308 16458
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13372 13938 13400 14214
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12707 13084 13015 13093
rect 12707 13082 12713 13084
rect 12769 13082 12793 13084
rect 12849 13082 12873 13084
rect 12929 13082 12953 13084
rect 13009 13082 13015 13084
rect 12769 13030 12771 13082
rect 12951 13030 12953 13082
rect 12707 13028 12713 13030
rect 12769 13028 12793 13030
rect 12849 13028 12873 13030
rect 12929 13028 12953 13030
rect 13009 13028 13015 13030
rect 12707 13019 13015 13028
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12636 12838 12756 12866
rect 12728 12434 12756 12838
rect 12820 12753 12848 12922
rect 12806 12744 12862 12753
rect 12806 12679 12862 12688
rect 13096 12481 13124 13518
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13082 12472 13138 12481
rect 12452 12406 12572 12434
rect 12728 12406 13032 12434
rect 13082 12407 13138 12416
rect 12438 12336 12494 12345
rect 12438 12271 12494 12280
rect 12452 11937 12480 12271
rect 12438 11928 12494 11937
rect 12438 11863 12494 11872
rect 12438 11520 12494 11529
rect 12047 11452 12355 11461
rect 12438 11455 12494 11464
rect 12047 11450 12053 11452
rect 12109 11450 12133 11452
rect 12189 11450 12213 11452
rect 12269 11450 12293 11452
rect 12349 11450 12355 11452
rect 12109 11398 12111 11450
rect 12291 11398 12293 11450
rect 12047 11396 12053 11398
rect 12109 11396 12133 11398
rect 12189 11396 12213 11398
rect 12269 11396 12293 11398
rect 12349 11396 12355 11398
rect 12047 11387 12355 11396
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 12176 10606 12204 11086
rect 12452 10849 12480 11455
rect 12438 10840 12494 10849
rect 12438 10775 12494 10784
rect 12438 10704 12494 10713
rect 12438 10639 12494 10648
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11992 10418 12020 10542
rect 12452 10441 12480 10639
rect 11900 10390 12020 10418
rect 12438 10432 12494 10441
rect 11900 9738 11928 10390
rect 12047 10364 12355 10373
rect 12438 10367 12494 10376
rect 12047 10362 12053 10364
rect 12109 10362 12133 10364
rect 12189 10362 12213 10364
rect 12269 10362 12293 10364
rect 12349 10362 12355 10364
rect 12109 10310 12111 10362
rect 12291 10310 12293 10362
rect 12047 10308 12053 10310
rect 12109 10308 12133 10310
rect 12189 10308 12213 10310
rect 12269 10308 12293 10310
rect 12349 10308 12355 10310
rect 12047 10299 12355 10308
rect 12438 10296 12494 10305
rect 11980 10260 12032 10266
rect 12438 10231 12494 10240
rect 11980 10202 12032 10208
rect 11992 10062 12020 10202
rect 12452 10146 12480 10231
rect 12176 10130 12480 10146
rect 12164 10124 12480 10130
rect 12216 10118 12480 10124
rect 12164 10066 12216 10072
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 11900 9710 12020 9738
rect 11796 9648 11848 9654
rect 11702 9616 11758 9625
rect 11612 9580 11664 9586
rect 11796 9590 11848 9596
rect 11886 9616 11942 9625
rect 11702 9551 11758 9560
rect 11886 9551 11942 9560
rect 11612 9522 11664 9528
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 7750 11560 9046
rect 11624 8974 11652 9522
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11612 8832 11664 8838
rect 11610 8800 11612 8809
rect 11664 8800 11666 8809
rect 11610 8735 11666 8744
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11624 7750 11652 8570
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11518 7576 11574 7585
rect 11518 7511 11574 7520
rect 11532 7274 11560 7511
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11532 6322 11560 7210
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11624 3942 11652 7686
rect 11716 7002 11744 9551
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11808 9217 11836 9318
rect 11794 9208 11850 9217
rect 11794 9143 11850 9152
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11808 8566 11836 8842
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 11164 3466 11192 3674
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 10690 3088 10746 3097
rect 10796 3058 10824 3402
rect 10690 3023 10692 3032
rect 10744 3023 10746 3032
rect 10784 3052 10836 3058
rect 10692 2994 10744 3000
rect 10784 2994 10836 3000
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 11072 2446 11100 2790
rect 11164 2650 11192 3402
rect 11612 2984 11664 2990
rect 11242 2952 11298 2961
rect 11612 2926 11664 2932
rect 11242 2887 11298 2896
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10324 2440 10376 2446
rect 11060 2440 11112 2446
rect 10324 2382 10376 2388
rect 10980 2388 11060 2394
rect 10980 2382 11112 2388
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 10336 800 10364 2382
rect 10980 2366 11100 2382
rect 10980 800 11008 2366
rect 11256 1970 11284 2887
rect 11244 1964 11296 1970
rect 11244 1906 11296 1912
rect 11624 800 11652 2926
rect 11716 2038 11744 5510
rect 11808 3602 11836 6666
rect 11900 6322 11928 9551
rect 11992 9382 12020 9710
rect 11980 9376 12032 9382
rect 12360 9364 12388 9862
rect 12544 9738 12572 12406
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12636 11150 12664 12242
rect 13004 12186 13032 12406
rect 13004 12158 13216 12186
rect 12707 11996 13015 12005
rect 12707 11994 12713 11996
rect 12769 11994 12793 11996
rect 12849 11994 12873 11996
rect 12929 11994 12953 11996
rect 13009 11994 13015 11996
rect 12769 11942 12771 11994
rect 12951 11942 12953 11994
rect 12707 11940 12713 11942
rect 12769 11940 12793 11942
rect 12849 11940 12873 11942
rect 12929 11940 12953 11942
rect 13009 11940 13015 11942
rect 12707 11931 13015 11940
rect 12898 11792 12954 11801
rect 12898 11727 12954 11736
rect 12912 11626 12940 11727
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12636 10810 12664 11086
rect 12707 10908 13015 10917
rect 12707 10906 12713 10908
rect 12769 10906 12793 10908
rect 12849 10906 12873 10908
rect 12929 10906 12953 10908
rect 13009 10906 13015 10908
rect 12769 10854 12771 10906
rect 12951 10854 12953 10906
rect 12707 10852 12713 10854
rect 12769 10852 12793 10854
rect 12849 10852 12873 10854
rect 12929 10852 12953 10854
rect 13009 10852 13015 10854
rect 12707 10843 13015 10852
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12452 9710 12572 9738
rect 12452 9625 12480 9710
rect 12636 9674 12664 10474
rect 12820 10169 12848 10610
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13004 10169 13032 10542
rect 12806 10160 12862 10169
rect 12806 10095 12862 10104
rect 12990 10160 13046 10169
rect 12990 10095 13046 10104
rect 13096 9908 13124 11630
rect 13188 10062 13216 12158
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13280 10849 13308 12106
rect 13372 11529 13400 13874
rect 13464 13326 13492 16934
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13556 16114 13584 16390
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13556 14074 13584 16050
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13648 13954 13676 16934
rect 13832 16726 13860 17614
rect 14370 17575 14426 17584
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14292 15473 14320 16050
rect 14278 15464 14334 15473
rect 14278 15399 14334 15408
rect 14096 15360 14148 15366
rect 14280 15360 14332 15366
rect 14148 15308 14228 15314
rect 14096 15302 14228 15308
rect 14280 15302 14332 15308
rect 14108 15286 14228 15302
rect 14200 15026 14228 15286
rect 14292 15094 14320 15302
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14094 14920 14150 14929
rect 14094 14855 14150 14864
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13556 13926 13676 13954
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13556 13258 13584 13926
rect 13636 13864 13688 13870
rect 13740 13841 13768 14758
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13832 14278 13860 14350
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13636 13806 13688 13812
rect 13726 13832 13782 13841
rect 13648 13530 13676 13806
rect 13726 13767 13782 13776
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13740 13530 13768 13670
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13464 11937 13492 13126
rect 13556 12764 13584 13194
rect 13648 12918 13676 13466
rect 13740 12986 13768 13466
rect 13832 13433 13860 14214
rect 13924 13870 13952 14486
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13818 13424 13874 13433
rect 13818 13359 13874 13368
rect 13924 13161 13952 13466
rect 13910 13152 13966 13161
rect 13910 13087 13966 13096
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 14016 12850 14044 14010
rect 14108 14006 14136 14855
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14108 13258 14136 13942
rect 14200 13705 14228 14962
rect 14384 14618 14412 17575
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15212 16674 15240 17206
rect 15212 16658 15332 16674
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 15200 16652 15332 16658
rect 15252 16646 15332 16652
rect 15200 16594 15252 16600
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14568 15337 14596 16390
rect 14648 15360 14700 15366
rect 14554 15328 14610 15337
rect 14648 15302 14700 15308
rect 14554 15263 14610 15272
rect 14660 14906 14688 15302
rect 14568 14878 14688 14906
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14292 13802 14320 14282
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14186 13696 14242 13705
rect 14186 13631 14242 13640
rect 14292 13376 14320 13738
rect 14200 13348 14320 13376
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14094 13152 14150 13161
rect 14094 13087 14150 13096
rect 14108 12866 14136 13087
rect 14200 12986 14228 13348
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14004 12844 14056 12850
rect 14108 12838 14228 12866
rect 14004 12786 14056 12792
rect 13912 12776 13964 12782
rect 13556 12736 13768 12764
rect 13544 12640 13596 12646
rect 13740 12617 13768 12736
rect 13912 12718 13964 12724
rect 13820 12640 13872 12646
rect 13544 12582 13596 12588
rect 13726 12608 13782 12617
rect 13450 11928 13506 11937
rect 13450 11863 13506 11872
rect 13358 11520 13414 11529
rect 13358 11455 13414 11464
rect 13358 11112 13414 11121
rect 13358 11047 13414 11056
rect 13452 11076 13504 11082
rect 13266 10840 13322 10849
rect 13266 10775 13322 10784
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13268 9920 13320 9926
rect 13096 9880 13216 9908
rect 12707 9820 13015 9829
rect 12707 9818 12713 9820
rect 12769 9818 12793 9820
rect 12849 9818 12873 9820
rect 12929 9818 12953 9820
rect 13009 9818 13015 9820
rect 12769 9766 12771 9818
rect 12951 9766 12953 9818
rect 12707 9764 12713 9766
rect 12769 9764 12793 9766
rect 12849 9764 12873 9766
rect 12929 9764 12953 9766
rect 13009 9764 13015 9766
rect 12707 9755 13015 9764
rect 12636 9646 12848 9674
rect 12438 9616 12494 9625
rect 12438 9551 12494 9560
rect 12360 9336 12480 9364
rect 11980 9318 12032 9324
rect 12047 9276 12355 9285
rect 12047 9274 12053 9276
rect 12109 9274 12133 9276
rect 12189 9274 12213 9276
rect 12269 9274 12293 9276
rect 12349 9274 12355 9276
rect 12109 9222 12111 9274
rect 12291 9222 12293 9274
rect 12047 9220 12053 9222
rect 12109 9220 12133 9222
rect 12189 9220 12213 9222
rect 12269 9220 12293 9222
rect 12349 9220 12355 9222
rect 12047 9211 12355 9220
rect 12452 9160 12480 9336
rect 11992 9132 12480 9160
rect 12622 9208 12678 9217
rect 12622 9143 12678 9152
rect 11992 8294 12020 9132
rect 12636 8974 12664 9143
rect 12820 9024 12848 9646
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13004 9489 13032 9590
rect 12990 9480 13046 9489
rect 12990 9415 13046 9424
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12992 9036 13044 9042
rect 12820 8996 12992 9024
rect 12992 8978 13044 8984
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12624 8832 12676 8838
rect 12452 8792 12624 8820
rect 12452 8634 12480 8792
rect 12624 8774 12676 8780
rect 12707 8732 13015 8741
rect 12707 8730 12713 8732
rect 12769 8730 12793 8732
rect 12849 8730 12873 8732
rect 12929 8730 12953 8732
rect 13009 8730 13015 8732
rect 12769 8678 12771 8730
rect 12951 8678 12953 8730
rect 12707 8676 12713 8678
rect 12769 8676 12793 8678
rect 12849 8676 12873 8678
rect 12929 8676 12953 8678
rect 13009 8676 13015 8678
rect 12530 8664 12586 8673
rect 12707 8667 13015 8676
rect 12440 8628 12492 8634
rect 12586 8608 12940 8616
rect 12530 8599 12940 8608
rect 12544 8588 12940 8599
rect 12440 8570 12492 8576
rect 12452 8480 12480 8570
rect 12406 8452 12480 8480
rect 12544 8486 12848 8514
rect 12912 8498 12940 8588
rect 12406 8378 12434 8452
rect 12544 8430 12572 8486
rect 12532 8424 12584 8430
rect 12406 8350 12480 8378
rect 12532 8366 12584 8372
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 12047 8188 12355 8197
rect 12047 8186 12053 8188
rect 12109 8186 12133 8188
rect 12189 8186 12213 8188
rect 12269 8186 12293 8188
rect 12349 8186 12355 8188
rect 12109 8134 12111 8186
rect 12291 8134 12293 8186
rect 12047 8132 12053 8134
rect 12109 8132 12133 8134
rect 12189 8132 12213 8134
rect 12269 8132 12293 8134
rect 12349 8132 12355 8134
rect 12047 8123 12355 8132
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11992 7274 12020 7822
rect 12084 7274 12112 8026
rect 12268 7993 12296 8026
rect 12452 8004 12480 8350
rect 12530 8120 12586 8129
rect 12530 8055 12532 8064
rect 12584 8055 12586 8064
rect 12532 8026 12584 8032
rect 12254 7984 12310 7993
rect 12254 7919 12310 7928
rect 12406 7976 12480 8004
rect 12530 7984 12586 7993
rect 12406 7936 12434 7976
rect 12406 7908 12480 7936
rect 12530 7919 12586 7928
rect 12254 7848 12310 7857
rect 12254 7783 12310 7792
rect 12268 7750 12296 7783
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12162 7576 12218 7585
rect 12162 7511 12218 7520
rect 12176 7410 12204 7511
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 11980 7268 12032 7274
rect 11980 7210 12032 7216
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 6730 12204 6938
rect 12452 6905 12480 7908
rect 12544 7721 12572 7919
rect 12530 7712 12586 7721
rect 12530 7647 12586 7656
rect 12636 7546 12664 8366
rect 12820 8294 12848 8486
rect 12900 8492 12952 8498
rect 13096 8480 13124 9318
rect 13188 9092 13216 9880
rect 13268 9862 13320 9868
rect 13280 9722 13308 9862
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13280 9160 13308 9454
rect 13372 9353 13400 11047
rect 13452 11018 13504 11024
rect 13464 10606 13492 11018
rect 13556 10962 13584 12582
rect 13820 12582 13872 12588
rect 13726 12543 13782 12552
rect 13740 11762 13768 12543
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11150 13676 11494
rect 13726 11384 13782 11393
rect 13726 11319 13782 11328
rect 13740 11218 13768 11319
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13636 11144 13688 11150
rect 13832 11121 13860 12582
rect 13924 12442 13952 12718
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13924 11898 13952 12242
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13636 11086 13688 11092
rect 13818 11112 13874 11121
rect 13728 11076 13780 11082
rect 13818 11047 13874 11056
rect 13728 11018 13780 11024
rect 13556 10934 13676 10962
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13556 10674 13584 10746
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 13464 9897 13492 9930
rect 13450 9888 13506 9897
rect 13450 9823 13506 9832
rect 13556 9674 13584 10610
rect 13464 9646 13584 9674
rect 13464 9500 13492 9646
rect 13648 9610 13676 10934
rect 13740 9674 13768 11018
rect 13924 11014 13952 11834
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13924 10266 13952 10950
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13740 9646 13860 9674
rect 13636 9604 13688 9610
rect 13636 9546 13688 9552
rect 13544 9512 13596 9518
rect 13464 9472 13544 9500
rect 13544 9454 13596 9460
rect 13358 9344 13414 9353
rect 13358 9279 13414 9288
rect 13556 9160 13584 9454
rect 13832 9364 13860 9646
rect 14016 9586 14044 12786
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14108 9722 14136 12310
rect 14200 12102 14228 12838
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11762 14228 12038
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14200 10305 14228 10474
rect 14186 10296 14242 10305
rect 14186 10231 14242 10240
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14094 9616 14150 9625
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 14004 9580 14056 9586
rect 14094 9551 14150 9560
rect 14004 9522 14056 9528
rect 13740 9336 13860 9364
rect 13280 9132 13492 9160
rect 13556 9132 13676 9160
rect 13188 9064 13400 9092
rect 13096 8452 13308 8480
rect 12900 8434 12952 8440
rect 12820 8266 13124 8294
rect 12714 8256 12770 8265
rect 12714 8191 12770 8200
rect 12728 7818 12756 8191
rect 12806 7848 12862 7857
rect 12716 7812 12768 7818
rect 12806 7783 12862 7792
rect 12716 7754 12768 7760
rect 12820 7750 12848 7783
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 13096 7698 13124 8266
rect 13174 7712 13230 7721
rect 13096 7670 13174 7698
rect 12707 7644 13015 7653
rect 13174 7647 13230 7656
rect 12707 7642 12713 7644
rect 12769 7642 12793 7644
rect 12849 7642 12873 7644
rect 12929 7642 12953 7644
rect 13009 7642 13015 7644
rect 12769 7590 12771 7642
rect 12951 7590 12953 7642
rect 12707 7588 12713 7590
rect 12769 7588 12793 7590
rect 12849 7588 12873 7590
rect 12929 7588 12953 7590
rect 13009 7588 13015 7590
rect 12707 7579 13015 7588
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12912 6934 12940 7210
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 12716 6928 12768 6934
rect 12254 6896 12310 6905
rect 12254 6831 12310 6840
rect 12438 6896 12494 6905
rect 12716 6870 12768 6876
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12438 6831 12494 6840
rect 12268 6730 12296 6831
rect 12452 6798 12480 6831
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12622 6760 12678 6769
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12360 6633 12388 6666
rect 12346 6624 12402 6633
rect 12346 6559 12402 6568
rect 12544 6497 12572 6734
rect 12622 6695 12678 6704
rect 12530 6488 12586 6497
rect 12530 6423 12586 6432
rect 12636 6390 12664 6695
rect 12728 6662 12756 6870
rect 13004 6798 13032 6938
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12707 6556 13015 6565
rect 12707 6554 12713 6556
rect 12769 6554 12793 6556
rect 12849 6554 12873 6556
rect 12929 6554 12953 6556
rect 13009 6554 13015 6556
rect 12769 6502 12771 6554
rect 12951 6502 12953 6554
rect 12707 6500 12713 6502
rect 12769 6500 12793 6502
rect 12849 6500 12873 6502
rect 12929 6500 12953 6502
rect 13009 6500 13015 6502
rect 12707 6491 13015 6500
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 13096 6322 13124 6394
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12072 6180 12124 6186
rect 11900 6140 12072 6168
rect 11900 5710 11928 6140
rect 12072 6122 12124 6128
rect 12544 6089 12572 6258
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12820 6089 12848 6190
rect 12530 6080 12586 6089
rect 12047 6012 12355 6021
rect 12530 6015 12586 6024
rect 12806 6080 12862 6089
rect 12806 6015 12862 6024
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 12348 3664 12400 3670
rect 12346 3632 12348 3641
rect 12400 3632 12402 3641
rect 11796 3596 11848 3602
rect 12346 3567 12402 3576
rect 11796 3538 11848 3544
rect 11808 3097 11836 3538
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 11794 3088 11850 3097
rect 12360 3058 12388 3334
rect 12544 3194 12572 5850
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12636 4078 12664 5782
rect 12820 5778 12848 6015
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 13004 5574 13032 6190
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12707 5468 13015 5477
rect 12707 5466 12713 5468
rect 12769 5466 12793 5468
rect 12849 5466 12873 5468
rect 12929 5466 12953 5468
rect 13009 5466 13015 5468
rect 12769 5414 12771 5466
rect 12951 5414 12953 5466
rect 12707 5412 12713 5414
rect 12769 5412 12793 5414
rect 12849 5412 12873 5414
rect 12929 5412 12953 5414
rect 13009 5412 13015 5414
rect 12707 5403 13015 5412
rect 13096 4554 13124 5714
rect 13188 4826 13216 7278
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 12707 4380 13015 4389
rect 12707 4378 12713 4380
rect 12769 4378 12793 4380
rect 12849 4378 12873 4380
rect 12929 4378 12953 4380
rect 13009 4378 13015 4380
rect 12769 4326 12771 4378
rect 12951 4326 12953 4378
rect 12707 4324 12713 4326
rect 12769 4324 12793 4326
rect 12849 4324 12873 4326
rect 12929 4324 12953 4326
rect 13009 4324 13015 4326
rect 12707 4315 13015 4324
rect 12898 4176 12954 4185
rect 12898 4111 12954 4120
rect 13084 4140 13136 4146
rect 12912 4078 12940 4111
rect 13084 4082 13136 4088
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12636 3194 12664 3470
rect 12707 3292 13015 3301
rect 12707 3290 12713 3292
rect 12769 3290 12793 3292
rect 12849 3290 12873 3292
rect 12929 3290 12953 3292
rect 13009 3290 13015 3292
rect 12769 3238 12771 3290
rect 12951 3238 12953 3290
rect 12707 3236 12713 3238
rect 12769 3236 12793 3238
rect 12849 3236 12873 3238
rect 12929 3236 12953 3238
rect 13009 3236 13015 3238
rect 12707 3227 13015 3236
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 11794 3023 11850 3032
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12360 2836 12388 2994
rect 13096 2990 13124 4082
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13188 3058 13216 3606
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 12360 2808 12480 2836
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 12452 2632 12480 2808
rect 12268 2604 12480 2632
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 12084 1902 12112 2314
rect 12072 1896 12124 1902
rect 12072 1838 12124 1844
rect 12268 800 12296 2604
rect 12636 2514 12664 2926
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12820 2310 12848 2450
rect 12808 2304 12860 2310
rect 13280 2292 13308 8452
rect 13372 7002 13400 9064
rect 13464 8945 13492 9132
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13450 8936 13506 8945
rect 13450 8871 13506 8880
rect 13556 8820 13584 8978
rect 13648 8974 13676 9132
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13464 8792 13584 8820
rect 13464 8090 13492 8792
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7410 13492 7686
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13464 7154 13492 7346
rect 13556 7274 13584 8298
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 13648 7206 13676 8366
rect 13740 7954 13768 9336
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13832 9081 13860 9114
rect 13818 9072 13874 9081
rect 13818 9007 13874 9016
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8401 13860 8910
rect 13818 8392 13874 8401
rect 13818 8327 13874 8336
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13726 7304 13782 7313
rect 13726 7239 13728 7248
rect 13780 7239 13782 7248
rect 13728 7210 13780 7216
rect 13636 7200 13688 7206
rect 13464 7126 13584 7154
rect 13636 7142 13688 7148
rect 13450 7032 13506 7041
rect 13360 6996 13412 7002
rect 13450 6967 13506 6976
rect 13360 6938 13412 6944
rect 13358 6896 13414 6905
rect 13358 6831 13414 6840
rect 13372 6798 13400 6831
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13372 3602 13400 3878
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13372 2650 13400 3130
rect 13464 2990 13492 6967
rect 13556 5914 13584 7126
rect 13648 6866 13676 7142
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13648 5778 13676 6802
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13648 3738 13676 4490
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13740 3602 13768 6870
rect 13832 6662 13860 8026
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13924 5574 13952 9522
rect 14108 9518 14136 9551
rect 14096 9512 14148 9518
rect 14002 9480 14058 9489
rect 14096 9454 14148 9460
rect 14002 9415 14058 9424
rect 14016 8809 14044 9415
rect 14200 8838 14228 10231
rect 14292 9194 14320 13194
rect 14384 11121 14412 14350
rect 14568 14006 14596 14878
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 12442 14504 13806
rect 14568 13161 14596 13942
rect 14554 13152 14610 13161
rect 14554 13087 14610 13096
rect 14464 12436 14516 12442
rect 14660 12434 14688 14758
rect 14752 13394 14780 16594
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15028 14890 15056 15302
rect 15304 15162 15332 16646
rect 15396 16250 15424 17983
rect 15566 17912 15622 17921
rect 15566 17847 15622 17856
rect 15580 16250 15608 17847
rect 17958 17776 18014 17785
rect 17958 17711 18014 17720
rect 17146 17436 17454 17445
rect 17146 17434 17152 17436
rect 17208 17434 17232 17436
rect 17288 17434 17312 17436
rect 17368 17434 17392 17436
rect 17448 17434 17454 17436
rect 17208 17382 17210 17434
rect 17390 17382 17392 17434
rect 17146 17380 17152 17382
rect 17208 17380 17232 17382
rect 17288 17380 17312 17382
rect 17368 17380 17392 17382
rect 17448 17380 17454 17382
rect 17146 17371 17454 17380
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16040 16794 16068 17070
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16316 16794 16344 16934
rect 16486 16892 16794 16901
rect 16486 16890 16492 16892
rect 16548 16890 16572 16892
rect 16628 16890 16652 16892
rect 16708 16890 16732 16892
rect 16788 16890 16794 16892
rect 16548 16838 16550 16890
rect 16730 16838 16732 16890
rect 16486 16836 16492 16838
rect 16548 16836 16572 16838
rect 16628 16836 16652 16838
rect 16708 16836 16732 16838
rect 16788 16836 16794 16838
rect 16486 16827 16794 16836
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 15750 16688 15806 16697
rect 15750 16623 15752 16632
rect 15804 16623 15806 16632
rect 15752 16594 15804 16600
rect 16040 16590 16068 16730
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15016 14884 15068 14890
rect 15016 14826 15068 14832
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 13870 14964 14758
rect 15028 13870 15056 14826
rect 15304 14822 15332 14962
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14936 13705 14964 13806
rect 14922 13696 14978 13705
rect 14922 13631 14978 13640
rect 15396 13530 15424 14486
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15212 13410 15240 13466
rect 15212 13394 15424 13410
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 15016 13388 15068 13394
rect 15212 13388 15436 13394
rect 15212 13382 15384 13388
rect 15016 13330 15068 13336
rect 15488 13376 15516 16118
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16028 15088 16080 15094
rect 16028 15030 16080 15036
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15566 14512 15622 14521
rect 15566 14447 15622 14456
rect 15580 14414 15608 14447
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15436 13348 15516 13376
rect 15384 13330 15436 13336
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14464 12378 14516 12384
rect 14568 12406 14688 12434
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11694 14504 12038
rect 14464 11688 14516 11694
rect 14462 11656 14464 11665
rect 14516 11656 14518 11665
rect 14462 11591 14518 11600
rect 14568 11234 14596 12406
rect 14844 12238 14872 12786
rect 14832 12232 14884 12238
rect 14936 12209 14964 13126
rect 15028 12782 15056 13330
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14832 12174 14884 12180
rect 14922 12200 14978 12209
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14476 11206 14596 11234
rect 14370 11112 14426 11121
rect 14370 11047 14426 11056
rect 14476 10554 14504 11206
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14568 10742 14596 11086
rect 14660 10742 14688 11086
rect 14752 10826 14780 11698
rect 14844 11014 14872 12174
rect 14922 12135 14978 12144
rect 15028 11354 15056 12718
rect 15120 12617 15148 12786
rect 15106 12608 15162 12617
rect 15106 12543 15162 12552
rect 15212 12050 15240 12854
rect 15304 12646 15332 13262
rect 15672 13138 15700 14214
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15396 13110 15700 13138
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15290 12472 15346 12481
rect 15290 12407 15346 12416
rect 15304 12102 15332 12407
rect 15120 12022 15240 12050
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15014 11248 15070 11257
rect 15014 11183 15070 11192
rect 14924 11144 14976 11150
rect 14922 11112 14924 11121
rect 14976 11112 14978 11121
rect 14922 11047 14978 11056
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14752 10798 14964 10826
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14738 10568 14794 10577
rect 14476 10526 14596 10554
rect 14462 10432 14518 10441
rect 14462 10367 14518 10376
rect 14476 9994 14504 10367
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14384 9489 14412 9658
rect 14370 9480 14426 9489
rect 14370 9415 14426 9424
rect 14372 9376 14424 9382
rect 14370 9344 14372 9353
rect 14424 9344 14426 9353
rect 14370 9279 14426 9288
rect 14292 9166 14412 9194
rect 14188 8832 14240 8838
rect 14002 8800 14058 8809
rect 14188 8774 14240 8780
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14002 8735 14058 8744
rect 14016 8634 14044 8735
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14188 8424 14240 8430
rect 14002 8392 14058 8401
rect 14188 8366 14240 8372
rect 14002 8327 14058 8336
rect 14016 6322 14044 8327
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7342 14136 7686
rect 14200 7546 14228 8366
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14002 5944 14058 5953
rect 14002 5879 14058 5888
rect 14016 5710 14044 5879
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14108 5642 14136 6734
rect 14186 6216 14242 6225
rect 14186 6151 14242 6160
rect 14200 5914 14228 6151
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 14108 4690 14136 5578
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13832 2378 13860 4218
rect 14108 3466 14136 4626
rect 14292 4078 14320 8774
rect 14384 8090 14412 9166
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14384 7546 14412 8026
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14384 4758 14412 7482
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14476 4622 14504 9930
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14568 3641 14596 10526
rect 14738 10503 14794 10512
rect 14752 10470 14780 10503
rect 14648 10464 14700 10470
rect 14646 10432 14648 10441
rect 14740 10464 14792 10470
rect 14700 10432 14702 10441
rect 14740 10406 14792 10412
rect 14646 10367 14702 10376
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14660 7970 14688 9998
rect 14752 8401 14780 10406
rect 14936 10130 14964 10798
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14844 9178 14872 10066
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14936 8838 14964 10066
rect 15028 8974 15056 11183
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15120 8906 15148 12022
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 9081 15240 10950
rect 15198 9072 15254 9081
rect 15198 9007 15254 9016
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14738 8392 14794 8401
rect 14738 8327 14794 8336
rect 14660 7942 14872 7970
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14752 7750 14780 7822
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14646 6896 14702 6905
rect 14646 6831 14702 6840
rect 14660 3670 14688 6831
rect 14752 6458 14780 7686
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14844 5030 14872 7942
rect 14936 7818 14964 8774
rect 15108 8288 15160 8294
rect 15014 8256 15070 8265
rect 15108 8230 15160 8236
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15014 8191 15070 8200
rect 15028 8022 15056 8191
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 15120 7818 15148 8230
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14844 4826 14872 4966
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14648 3664 14700 3670
rect 14554 3632 14610 3641
rect 14464 3596 14516 3602
rect 14648 3606 14700 3612
rect 14554 3567 14610 3576
rect 14464 3538 14516 3544
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 14108 2990 14136 3402
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14004 2644 14056 2650
rect 14372 2644 14424 2650
rect 14056 2604 14372 2632
rect 14004 2586 14056 2592
rect 14372 2586 14424 2592
rect 14476 2582 14504 3538
rect 14464 2576 14516 2582
rect 14464 2518 14516 2524
rect 14568 2446 14596 3567
rect 14936 3126 14964 7754
rect 15106 7712 15162 7721
rect 15106 7647 15162 7656
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15028 3738 15056 7346
rect 15120 5642 15148 7647
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 4214 15148 5578
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 15212 3738 15240 8230
rect 15304 4146 15332 11290
rect 15396 9382 15424 13110
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15488 12170 15516 12922
rect 15566 12744 15622 12753
rect 15566 12679 15568 12688
rect 15620 12679 15622 12688
rect 15568 12650 15620 12656
rect 15764 12646 15792 13330
rect 15856 12986 15884 14214
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15752 12640 15804 12646
rect 15566 12608 15622 12617
rect 15752 12582 15804 12588
rect 15566 12543 15622 12552
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15488 11801 15516 11834
rect 15474 11792 15530 11801
rect 15474 11727 15530 11736
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15396 8566 15424 9114
rect 15488 8906 15516 11727
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15304 3194 15332 4082
rect 15396 4049 15424 8298
rect 15580 8242 15608 12543
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15672 12238 15700 12378
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15672 11801 15700 12174
rect 15658 11792 15714 11801
rect 15658 11727 15714 11736
rect 15764 11082 15792 12582
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15672 9178 15700 9454
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15658 8936 15714 8945
rect 15658 8871 15714 8880
rect 15488 8214 15608 8242
rect 15488 7546 15516 8214
rect 15566 8120 15622 8129
rect 15566 8055 15622 8064
rect 15580 7954 15608 8055
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15580 7002 15608 7754
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15474 5672 15530 5681
rect 15474 5607 15530 5616
rect 15488 4146 15516 5607
rect 15672 5302 15700 8871
rect 15764 8090 15792 10202
rect 15856 8634 15884 12786
rect 15948 12628 15976 14758
rect 16040 14362 16068 15030
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16132 14482 16160 14894
rect 16224 14482 16252 15098
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16040 14334 16160 14362
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16040 12850 16068 13466
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15948 12600 16068 12628
rect 15934 12336 15990 12345
rect 15934 12271 15936 12280
rect 15988 12271 15990 12280
rect 15936 12242 15988 12248
rect 15948 11354 15976 12242
rect 16040 11558 16068 12600
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16040 11286 16068 11494
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16132 11098 16160 14334
rect 16224 14074 16252 14418
rect 16316 14346 16344 16730
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16684 16250 16712 16526
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16486 15804 16794 15813
rect 16486 15802 16492 15804
rect 16548 15802 16572 15804
rect 16628 15802 16652 15804
rect 16708 15802 16732 15804
rect 16788 15802 16794 15804
rect 16548 15750 16550 15802
rect 16730 15750 16732 15802
rect 16486 15748 16492 15750
rect 16548 15748 16572 15750
rect 16628 15748 16652 15750
rect 16708 15748 16732 15750
rect 16788 15748 16794 15750
rect 16486 15739 16794 15748
rect 16868 15570 16896 16390
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 16304 14340 16356 14346
rect 16304 14282 16356 14288
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16224 12782 16252 14010
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16316 12434 16344 13806
rect 16408 12986 16436 15370
rect 16486 14716 16794 14725
rect 16486 14714 16492 14716
rect 16548 14714 16572 14716
rect 16628 14714 16652 14716
rect 16708 14714 16732 14716
rect 16788 14714 16794 14716
rect 16548 14662 16550 14714
rect 16730 14662 16732 14714
rect 16486 14660 16492 14662
rect 16548 14660 16572 14662
rect 16628 14660 16652 14662
rect 16708 14660 16732 14662
rect 16788 14660 16794 14662
rect 16486 14651 16794 14660
rect 16486 13628 16794 13637
rect 16486 13626 16492 13628
rect 16548 13626 16572 13628
rect 16628 13626 16652 13628
rect 16708 13626 16732 13628
rect 16788 13626 16794 13628
rect 16548 13574 16550 13626
rect 16730 13574 16732 13626
rect 16486 13572 16492 13574
rect 16548 13572 16572 13574
rect 16628 13572 16652 13574
rect 16708 13572 16732 13574
rect 16788 13572 16794 13574
rect 16486 13563 16794 13572
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16396 12776 16448 12782
rect 16500 12753 16528 13262
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16684 12850 16712 13194
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16396 12718 16448 12724
rect 16486 12744 16542 12753
rect 15948 11070 16160 11098
rect 16224 12406 16344 12434
rect 15948 10146 15976 11070
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16040 10266 16068 10406
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15948 10118 16068 10146
rect 16040 9722 16068 10118
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16026 9480 16082 9489
rect 15936 9444 15988 9450
rect 16026 9415 16082 9424
rect 15936 9386 15988 9392
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15764 7478 15792 8026
rect 15856 7750 15884 8230
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15382 4040 15438 4049
rect 15382 3975 15438 3984
rect 15488 3890 15516 4082
rect 15488 3862 15608 3890
rect 15474 3768 15530 3777
rect 15474 3703 15476 3712
rect 15528 3703 15530 3712
rect 15476 3674 15528 3680
rect 15580 3466 15608 3862
rect 15856 3602 15884 7482
rect 15948 6934 15976 9386
rect 16040 9178 16068 9415
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 16040 8430 16068 8842
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16040 8090 16068 8366
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16040 7546 16068 8026
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 16040 6186 16068 7278
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 16132 4554 16160 10950
rect 16224 10470 16252 12406
rect 16408 11898 16436 12718
rect 16960 12696 16988 17274
rect 17774 16552 17830 16561
rect 17774 16487 17830 16496
rect 17146 16348 17454 16357
rect 17146 16346 17152 16348
rect 17208 16346 17232 16348
rect 17288 16346 17312 16348
rect 17368 16346 17392 16348
rect 17448 16346 17454 16348
rect 17208 16294 17210 16346
rect 17390 16294 17392 16346
rect 17146 16292 17152 16294
rect 17208 16292 17232 16294
rect 17288 16292 17312 16294
rect 17368 16292 17392 16294
rect 17448 16292 17454 16294
rect 17146 16283 17454 16292
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17146 15260 17454 15269
rect 17146 15258 17152 15260
rect 17208 15258 17232 15260
rect 17288 15258 17312 15260
rect 17368 15258 17392 15260
rect 17448 15258 17454 15260
rect 17208 15206 17210 15258
rect 17390 15206 17392 15258
rect 17146 15204 17152 15206
rect 17208 15204 17232 15206
rect 17288 15204 17312 15206
rect 17368 15204 17392 15206
rect 17448 15204 17454 15206
rect 17146 15195 17454 15204
rect 17498 14376 17554 14385
rect 17498 14311 17554 14320
rect 17146 14172 17454 14181
rect 17146 14170 17152 14172
rect 17208 14170 17232 14172
rect 17288 14170 17312 14172
rect 17368 14170 17392 14172
rect 17448 14170 17454 14172
rect 17208 14118 17210 14170
rect 17390 14118 17392 14170
rect 17146 14116 17152 14118
rect 17208 14116 17232 14118
rect 17288 14116 17312 14118
rect 17368 14116 17392 14118
rect 17448 14116 17454 14118
rect 17146 14107 17454 14116
rect 17146 13084 17454 13093
rect 17146 13082 17152 13084
rect 17208 13082 17232 13084
rect 17288 13082 17312 13084
rect 17368 13082 17392 13084
rect 17448 13082 17454 13084
rect 17208 13030 17210 13082
rect 17390 13030 17392 13082
rect 17146 13028 17152 13030
rect 17208 13028 17232 13030
rect 17288 13028 17312 13030
rect 17368 13028 17392 13030
rect 17448 13028 17454 13030
rect 17146 13019 17454 13028
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 16486 12679 16542 12688
rect 16868 12668 16988 12696
rect 16486 12540 16794 12549
rect 16486 12538 16492 12540
rect 16548 12538 16572 12540
rect 16628 12538 16652 12540
rect 16708 12538 16732 12540
rect 16788 12538 16794 12540
rect 16548 12486 16550 12538
rect 16730 12486 16732 12538
rect 16486 12484 16492 12486
rect 16548 12484 16572 12486
rect 16628 12484 16652 12486
rect 16708 12484 16732 12486
rect 16788 12484 16794 12486
rect 16486 12475 16794 12484
rect 16868 11898 16896 12668
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16304 11824 16356 11830
rect 16488 11824 16540 11830
rect 16304 11766 16356 11772
rect 16394 11792 16450 11801
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 9926 16252 10406
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16224 9382 16252 9658
rect 16316 9654 16344 11766
rect 16450 11772 16488 11778
rect 16450 11766 16540 11772
rect 16450 11750 16528 11766
rect 16948 11756 17000 11762
rect 16394 11727 16450 11736
rect 16408 11336 16436 11727
rect 16948 11698 17000 11704
rect 16486 11452 16794 11461
rect 16486 11450 16492 11452
rect 16548 11450 16572 11452
rect 16628 11450 16652 11452
rect 16708 11450 16732 11452
rect 16788 11450 16794 11452
rect 16548 11398 16550 11450
rect 16730 11398 16732 11450
rect 16486 11396 16492 11398
rect 16548 11396 16572 11398
rect 16628 11396 16652 11398
rect 16708 11396 16732 11398
rect 16788 11396 16794 11398
rect 16486 11387 16794 11396
rect 16408 11308 16528 11336
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16408 10577 16436 11086
rect 16500 10674 16528 11308
rect 16672 11280 16724 11286
rect 16960 11257 16988 11698
rect 16672 11222 16724 11228
rect 16946 11248 17002 11257
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16592 10713 16620 11086
rect 16578 10704 16634 10713
rect 16488 10668 16540 10674
rect 16684 10674 16712 11222
rect 16946 11183 17002 11192
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16854 10976 16910 10985
rect 16854 10911 16910 10920
rect 16762 10840 16818 10849
rect 16762 10775 16764 10784
rect 16816 10775 16818 10784
rect 16764 10746 16816 10752
rect 16578 10639 16634 10648
rect 16672 10668 16724 10674
rect 16488 10610 16540 10616
rect 16672 10610 16724 10616
rect 16394 10568 16450 10577
rect 16394 10503 16450 10512
rect 16500 10452 16528 10610
rect 16408 10424 16528 10452
rect 16408 10062 16436 10424
rect 16486 10364 16794 10373
rect 16486 10362 16492 10364
rect 16548 10362 16572 10364
rect 16628 10362 16652 10364
rect 16708 10362 16732 10364
rect 16788 10362 16794 10364
rect 16548 10310 16550 10362
rect 16730 10310 16732 10362
rect 16486 10308 16492 10310
rect 16548 10308 16572 10310
rect 16628 10308 16652 10310
rect 16708 10308 16732 10310
rect 16788 10308 16794 10310
rect 16486 10299 16794 10308
rect 16868 10146 16896 10911
rect 16776 10118 16896 10146
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 5681 16252 9318
rect 16316 8974 16344 9454
rect 16408 9110 16436 9998
rect 16486 9616 16542 9625
rect 16486 9551 16542 9560
rect 16500 9518 16528 9551
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16776 9382 16804 10118
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16868 9568 16896 9930
rect 16960 9761 16988 11086
rect 17052 10538 17080 12922
rect 17222 12880 17278 12889
rect 17512 12850 17540 14311
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17222 12815 17224 12824
rect 17276 12815 17278 12824
rect 17500 12844 17552 12850
rect 17224 12786 17276 12792
rect 17500 12786 17552 12792
rect 17146 11996 17454 12005
rect 17146 11994 17152 11996
rect 17208 11994 17232 11996
rect 17288 11994 17312 11996
rect 17368 11994 17392 11996
rect 17448 11994 17454 11996
rect 17208 11942 17210 11994
rect 17390 11942 17392 11994
rect 17146 11940 17152 11942
rect 17208 11940 17232 11942
rect 17288 11940 17312 11942
rect 17368 11940 17392 11942
rect 17448 11940 17454 11942
rect 17146 11931 17454 11940
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17328 11082 17356 11766
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17146 10908 17454 10917
rect 17146 10906 17152 10908
rect 17208 10906 17232 10908
rect 17288 10906 17312 10908
rect 17368 10906 17392 10908
rect 17448 10906 17454 10908
rect 17208 10854 17210 10906
rect 17390 10854 17392 10906
rect 17146 10852 17152 10854
rect 17208 10852 17232 10854
rect 17288 10852 17312 10854
rect 17368 10852 17392 10854
rect 17448 10852 17454 10854
rect 17146 10843 17454 10852
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17040 10532 17092 10538
rect 17040 10474 17092 10480
rect 17420 10062 17448 10610
rect 17408 10056 17460 10062
rect 17038 10024 17094 10033
rect 17408 9998 17460 10004
rect 17038 9959 17094 9968
rect 16946 9752 17002 9761
rect 16946 9687 17002 9696
rect 17052 9674 17080 9959
rect 17146 9820 17454 9829
rect 17146 9818 17152 9820
rect 17208 9818 17232 9820
rect 17288 9818 17312 9820
rect 17368 9818 17392 9820
rect 17448 9818 17454 9820
rect 17208 9766 17210 9818
rect 17390 9766 17392 9818
rect 17146 9764 17152 9766
rect 17208 9764 17232 9766
rect 17288 9764 17312 9766
rect 17368 9764 17392 9766
rect 17448 9764 17454 9766
rect 17146 9755 17454 9764
rect 17052 9646 17448 9674
rect 16844 9540 16896 9568
rect 16948 9580 17000 9586
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16486 9276 16794 9285
rect 16486 9274 16492 9276
rect 16548 9274 16572 9276
rect 16628 9274 16652 9276
rect 16708 9274 16732 9276
rect 16788 9274 16794 9276
rect 16548 9222 16550 9274
rect 16730 9222 16732 9274
rect 16486 9220 16492 9222
rect 16548 9220 16572 9222
rect 16628 9220 16652 9222
rect 16708 9220 16732 9222
rect 16788 9220 16794 9222
rect 16486 9211 16794 9220
rect 16396 9104 16448 9110
rect 16844 9092 16872 9540
rect 16948 9522 17000 9528
rect 16960 9489 16988 9522
rect 17316 9512 17368 9518
rect 16946 9480 17002 9489
rect 17316 9454 17368 9460
rect 16946 9415 17002 9424
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17052 9160 17080 9318
rect 16960 9132 17080 9160
rect 16844 9064 16896 9092
rect 16396 9046 16448 9052
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16316 7478 16344 8774
rect 16408 8430 16436 8910
rect 16776 8498 16804 8978
rect 16868 8634 16896 9064
rect 16960 8634 16988 9132
rect 17144 9024 17172 9318
rect 17328 9178 17356 9454
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17144 8996 17356 9024
rect 17328 8945 17356 8996
rect 17314 8936 17370 8945
rect 17040 8900 17092 8906
rect 17314 8871 17370 8880
rect 17040 8842 17092 8848
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16396 8424 16448 8430
rect 16948 8424 17000 8430
rect 16396 8366 16448 8372
rect 16854 8392 16910 8401
rect 16948 8366 17000 8372
rect 16854 8327 16910 8336
rect 16486 8188 16794 8197
rect 16486 8186 16492 8188
rect 16548 8186 16572 8188
rect 16628 8186 16652 8188
rect 16708 8186 16732 8188
rect 16788 8186 16794 8188
rect 16548 8134 16550 8186
rect 16730 8134 16732 8186
rect 16486 8132 16492 8134
rect 16548 8132 16572 8134
rect 16628 8132 16652 8134
rect 16708 8132 16732 8134
rect 16788 8132 16794 8134
rect 16486 8123 16794 8132
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16408 7721 16436 8026
rect 16868 7818 16896 8327
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16394 7712 16450 7721
rect 16960 7698 16988 8366
rect 17052 8090 17080 8842
rect 17420 8838 17448 9646
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17146 8732 17454 8741
rect 17146 8730 17152 8732
rect 17208 8730 17232 8732
rect 17288 8730 17312 8732
rect 17368 8730 17392 8732
rect 17448 8730 17454 8732
rect 17208 8678 17210 8730
rect 17390 8678 17392 8730
rect 17146 8676 17152 8678
rect 17208 8676 17232 8678
rect 17288 8676 17312 8678
rect 17368 8676 17392 8678
rect 17448 8676 17454 8678
rect 17146 8667 17454 8676
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17038 7984 17094 7993
rect 17038 7919 17094 7928
rect 16394 7647 16450 7656
rect 16868 7670 16988 7698
rect 16394 7576 16450 7585
rect 16394 7511 16450 7520
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16210 5672 16266 5681
rect 16210 5607 16266 5616
rect 16210 5264 16266 5273
rect 16210 5199 16266 5208
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15856 3194 15884 3538
rect 16224 3534 16252 5199
rect 16316 5166 16344 6938
rect 16408 6866 16436 7511
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 16868 6882 16896 7670
rect 17052 7546 17080 7919
rect 17144 7750 17172 8570
rect 17236 8498 17264 8570
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17512 8430 17540 11562
rect 17604 10742 17632 13126
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17590 10160 17646 10169
rect 17590 10095 17646 10104
rect 17316 8424 17368 8430
rect 17500 8424 17552 8430
rect 17316 8366 17368 8372
rect 17498 8392 17500 8401
rect 17552 8392 17554 8401
rect 17328 8022 17356 8366
rect 17498 8327 17554 8336
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17146 7644 17454 7653
rect 17146 7642 17152 7644
rect 17208 7642 17232 7644
rect 17288 7642 17312 7644
rect 17368 7642 17392 7644
rect 17448 7642 17454 7644
rect 17208 7590 17210 7642
rect 17390 7590 17392 7642
rect 17146 7588 17152 7590
rect 17208 7588 17232 7590
rect 17288 7588 17312 7590
rect 17368 7588 17392 7590
rect 17448 7588 17454 7590
rect 17146 7579 17454 7588
rect 17512 7546 17540 7822
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17038 7440 17094 7449
rect 17604 7426 17632 10095
rect 17696 8634 17724 15982
rect 17788 15502 17816 16487
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17788 15162 17816 15438
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17788 14113 17816 15098
rect 17880 14929 17908 15438
rect 17866 14920 17922 14929
rect 17866 14855 17922 14864
rect 17774 14104 17830 14113
rect 17774 14039 17830 14048
rect 17880 11286 17908 14855
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17774 9616 17830 9625
rect 17880 9602 17908 11018
rect 17972 10674 18000 17711
rect 18972 17604 19024 17610
rect 18972 17546 19024 17552
rect 18786 15600 18842 15609
rect 18786 15535 18842 15544
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18050 13288 18106 13297
rect 18050 13223 18106 13232
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9722 18000 9998
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17880 9574 18000 9602
rect 17774 9551 17830 9560
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17788 8498 17816 9551
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17094 7410 17172 7426
rect 17094 7404 17184 7410
rect 17094 7398 17132 7404
rect 17038 7375 17094 7384
rect 16396 6860 16448 6866
rect 16868 6854 16988 6882
rect 16396 6802 16448 6808
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 16868 5914 16896 6666
rect 16960 6662 16988 6854
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16960 6361 16988 6598
rect 17052 6458 17080 7375
rect 17132 7346 17184 7352
rect 17328 7398 17632 7426
rect 17328 7342 17356 7398
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17328 7002 17356 7278
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17316 6724 17368 6730
rect 17420 6712 17448 7278
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17368 6684 17448 6712
rect 17316 6666 17368 6672
rect 17146 6556 17454 6565
rect 17146 6554 17152 6556
rect 17208 6554 17232 6556
rect 17288 6554 17312 6556
rect 17368 6554 17392 6556
rect 17448 6554 17454 6556
rect 17208 6502 17210 6554
rect 17390 6502 17392 6554
rect 17146 6500 17152 6502
rect 17208 6500 17232 6502
rect 17288 6500 17312 6502
rect 17368 6500 17392 6502
rect 17448 6500 17454 6502
rect 17146 6491 17454 6500
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16946 6352 17002 6361
rect 16946 6287 17002 6296
rect 17498 6352 17554 6361
rect 17498 6287 17554 6296
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16394 5808 16450 5817
rect 16394 5743 16450 5752
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16408 4146 16436 5743
rect 17146 5468 17454 5477
rect 17146 5466 17152 5468
rect 17208 5466 17232 5468
rect 17288 5466 17312 5468
rect 17368 5466 17392 5468
rect 17448 5466 17454 5468
rect 17208 5414 17210 5466
rect 17390 5414 17392 5466
rect 17146 5412 17152 5414
rect 17208 5412 17232 5414
rect 17288 5412 17312 5414
rect 17368 5412 17392 5414
rect 17448 5412 17454 5414
rect 17146 5403 17454 5412
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 16854 4720 16910 4729
rect 16854 4655 16856 4664
rect 16908 4655 16910 4664
rect 16856 4626 16908 4632
rect 17512 4486 17540 6287
rect 17604 5914 17632 6802
rect 17696 6798 17724 8434
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17788 6458 17816 8298
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17880 6338 17908 9454
rect 17972 9042 18000 9574
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 18064 8514 18092 13223
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 17972 8498 18092 8514
rect 17960 8492 18092 8498
rect 18012 8486 18092 8492
rect 17960 8434 18012 8440
rect 17972 7478 18000 8434
rect 18050 7848 18106 7857
rect 18050 7783 18106 7792
rect 18064 7750 18092 7783
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17788 6310 17908 6338
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17788 5137 17816 6310
rect 17972 5370 18000 7278
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18064 5778 18092 6734
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17774 5128 17830 5137
rect 17774 5063 17830 5072
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17146 4380 17454 4389
rect 17146 4378 17152 4380
rect 17208 4378 17232 4380
rect 17288 4378 17312 4380
rect 17368 4378 17392 4380
rect 17448 4378 17454 4380
rect 17208 4326 17210 4378
rect 17390 4326 17392 4378
rect 17146 4324 17152 4326
rect 17208 4324 17232 4326
rect 17288 4324 17312 4326
rect 17368 4324 17392 4326
rect 17448 4324 17454 4326
rect 17146 4315 17454 4324
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16316 3602 16344 4014
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16408 3398 16436 3878
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 17420 3398 17448 4150
rect 17880 4146 17908 5034
rect 18064 5030 18092 5714
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18064 3602 18092 4966
rect 18156 4622 18184 11630
rect 18340 9602 18368 15302
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18616 12434 18644 13398
rect 18616 12406 18736 12434
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11150 18460 11494
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18432 10690 18460 11086
rect 18432 10674 18552 10690
rect 18420 10668 18552 10674
rect 18472 10662 18552 10668
rect 18420 10610 18472 10616
rect 18248 9574 18368 9602
rect 18420 9580 18472 9586
rect 18248 7750 18276 9574
rect 18420 9522 18472 9528
rect 18432 8634 18460 9522
rect 18524 9382 18552 10662
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18524 8514 18552 9318
rect 18602 9072 18658 9081
rect 18602 9007 18658 9016
rect 18432 8486 18552 8514
rect 18326 8392 18382 8401
rect 18326 8327 18382 8336
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15948 2922 15976 3334
rect 16408 3126 16436 3334
rect 17146 3292 17454 3301
rect 17146 3290 17152 3292
rect 17208 3290 17232 3292
rect 17288 3290 17312 3292
rect 17368 3290 17392 3292
rect 17448 3290 17454 3292
rect 17208 3238 17210 3290
rect 17390 3238 17392 3290
rect 17146 3236 17152 3238
rect 17208 3236 17232 3238
rect 17288 3236 17312 3238
rect 17368 3236 17392 3238
rect 17448 3236 17454 3238
rect 17146 3227 17454 3236
rect 17774 3224 17830 3233
rect 17774 3159 17776 3168
rect 17828 3159 17830 3168
rect 17776 3130 17828 3136
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 17314 3088 17370 3097
rect 17314 3023 17370 3032
rect 17328 2972 17356 3023
rect 17408 2984 17460 2990
rect 17328 2944 17408 2972
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 17328 2650 17356 2944
rect 17408 2926 17460 2932
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 18248 2582 18276 7482
rect 18340 5234 18368 8327
rect 18432 8022 18460 8486
rect 18512 8424 18564 8430
rect 18616 8412 18644 9007
rect 18564 8384 18644 8412
rect 18512 8366 18564 8372
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18432 7410 18460 7958
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18432 6118 18460 7346
rect 18524 6458 18552 8366
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18432 5234 18460 5850
rect 18708 5302 18736 12406
rect 18800 7342 18828 15535
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18892 5914 18920 10678
rect 18984 8294 19012 17546
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18432 3058 18460 5170
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18432 2774 18460 2994
rect 19076 2774 19104 14486
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19168 4758 19196 14350
rect 19260 7546 19288 15370
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19352 8537 19380 12854
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19338 8528 19394 8537
rect 19338 8463 19394 8472
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 19352 2990 19380 8463
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 18432 2746 18644 2774
rect 18616 2650 18644 2746
rect 18800 2746 19104 2774
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 18236 2576 18288 2582
rect 18236 2518 18288 2524
rect 14936 2446 14964 2518
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13360 2304 13412 2310
rect 13280 2264 13360 2292
rect 12808 2246 12860 2252
rect 13360 2246 13412 2252
rect 12707 2204 13015 2213
rect 12707 2202 12713 2204
rect 12769 2202 12793 2204
rect 12849 2202 12873 2204
rect 12929 2202 12953 2204
rect 13009 2202 13015 2204
rect 12769 2150 12771 2202
rect 12951 2150 12953 2202
rect 12707 2148 12713 2150
rect 12769 2148 12793 2150
rect 12849 2148 12873 2150
rect 12929 2148 12953 2150
rect 13009 2148 13015 2150
rect 12707 2139 13015 2148
rect 15120 2106 15148 2382
rect 18800 2378 18828 2746
rect 19444 2446 19472 10066
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 18788 2372 18840 2378
rect 18788 2314 18840 2320
rect 17146 2204 17454 2213
rect 17146 2202 17152 2204
rect 17208 2202 17232 2204
rect 17288 2202 17312 2204
rect 17368 2202 17392 2204
rect 17448 2202 17454 2204
rect 17208 2150 17210 2202
rect 17390 2150 17392 2202
rect 17146 2148 17152 2150
rect 17208 2148 17232 2150
rect 17288 2148 17312 2150
rect 17368 2148 17392 2150
rect 17448 2148 17454 2150
rect 17146 2139 17454 2148
rect 15108 2100 15160 2106
rect 15108 2042 15160 2048
rect 8496 734 8708 762
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
<< via2 >>
rect 2870 19080 2926 19136
rect 2778 18400 2834 18456
rect 938 17856 994 17912
rect 386 16632 442 16688
rect 938 16632 994 16688
rect 6734 18128 6790 18184
rect 2962 17720 3018 17776
rect 3835 17434 3891 17436
rect 3915 17434 3971 17436
rect 3995 17434 4051 17436
rect 4075 17434 4131 17436
rect 3835 17382 3881 17434
rect 3881 17382 3891 17434
rect 3915 17382 3945 17434
rect 3945 17382 3957 17434
rect 3957 17382 3971 17434
rect 3995 17382 4009 17434
rect 4009 17382 4021 17434
rect 4021 17382 4051 17434
rect 4075 17382 4085 17434
rect 4085 17382 4131 17434
rect 3835 17380 3891 17382
rect 3915 17380 3971 17382
rect 3995 17380 4051 17382
rect 4075 17380 4131 17382
rect 1490 16360 1546 16416
rect 846 15816 902 15872
rect 846 6024 902 6080
rect 846 4936 902 4992
rect 846 4256 902 4312
rect 846 3596 902 3632
rect 846 3576 848 3596
rect 848 3576 900 3596
rect 900 3576 902 3596
rect 846 2932 848 2952
rect 848 2932 900 2952
rect 900 2932 902 2952
rect 846 2896 902 2932
rect 1398 15000 1454 15056
rect 1214 14356 1216 14376
rect 1216 14356 1268 14376
rect 1268 14356 1270 14376
rect 1214 14320 1270 14356
rect 1398 13640 1454 13696
rect 1214 12824 1270 12880
rect 1398 12280 1454 12336
rect 1582 14320 1638 14376
rect 1582 13912 1638 13968
rect 2134 15952 2190 16008
rect 1214 12144 1270 12200
rect 1398 10920 1454 10976
rect 1398 10260 1454 10296
rect 1398 10240 1400 10260
rect 1400 10240 1452 10260
rect 1452 10240 1454 10260
rect 1582 12280 1638 12336
rect 1582 11600 1638 11656
rect 1582 10532 1638 10568
rect 1582 10512 1584 10532
rect 1584 10512 1636 10532
rect 1636 10512 1638 10532
rect 1490 9016 1546 9072
rect 1398 8916 1400 8936
rect 1400 8916 1452 8936
rect 1452 8916 1454 8936
rect 1398 8880 1454 8916
rect 1490 8608 1546 8664
rect 1030 4664 1086 4720
rect 1582 8200 1638 8256
rect 1582 6840 1638 6896
rect 1950 12960 2006 13016
rect 2410 15308 2412 15328
rect 2412 15308 2464 15328
rect 2464 15308 2466 15328
rect 2410 15272 2466 15308
rect 2778 16532 2780 16552
rect 2780 16532 2832 16552
rect 2832 16532 2834 16552
rect 2778 16496 2834 16532
rect 2778 16108 2834 16144
rect 2778 16088 2780 16108
rect 2780 16088 2832 16108
rect 2832 16088 2834 16108
rect 3054 17040 3110 17096
rect 2962 16496 3018 16552
rect 2502 15000 2558 15056
rect 2226 14456 2282 14512
rect 2686 14048 2742 14104
rect 2318 11192 2374 11248
rect 1950 9560 2006 9616
rect 1858 7404 1914 7440
rect 1858 7384 1860 7404
rect 1860 7384 1912 7404
rect 1912 7384 1914 7404
rect 1674 5752 1730 5808
rect 1582 5480 1638 5536
rect 2134 7520 2190 7576
rect 2134 7248 2190 7304
rect 3175 16890 3231 16892
rect 3255 16890 3311 16892
rect 3335 16890 3391 16892
rect 3415 16890 3471 16892
rect 3175 16838 3221 16890
rect 3221 16838 3231 16890
rect 3255 16838 3285 16890
rect 3285 16838 3297 16890
rect 3297 16838 3311 16890
rect 3335 16838 3349 16890
rect 3349 16838 3361 16890
rect 3361 16838 3391 16890
rect 3415 16838 3425 16890
rect 3425 16838 3471 16890
rect 3175 16836 3231 16838
rect 3255 16836 3311 16838
rect 3335 16836 3391 16838
rect 3415 16836 3471 16838
rect 3175 15802 3231 15804
rect 3255 15802 3311 15804
rect 3335 15802 3391 15804
rect 3415 15802 3471 15804
rect 3175 15750 3221 15802
rect 3221 15750 3231 15802
rect 3255 15750 3285 15802
rect 3285 15750 3297 15802
rect 3297 15750 3311 15802
rect 3335 15750 3349 15802
rect 3349 15750 3361 15802
rect 3361 15750 3391 15802
rect 3415 15750 3425 15802
rect 3425 15750 3471 15802
rect 3175 15748 3231 15750
rect 3255 15748 3311 15750
rect 3335 15748 3391 15750
rect 3415 15748 3471 15750
rect 5078 17040 5134 17096
rect 3882 16632 3938 16688
rect 3835 16346 3891 16348
rect 3915 16346 3971 16348
rect 3995 16346 4051 16348
rect 4075 16346 4131 16348
rect 3835 16294 3881 16346
rect 3881 16294 3891 16346
rect 3915 16294 3945 16346
rect 3945 16294 3957 16346
rect 3957 16294 3971 16346
rect 3995 16294 4009 16346
rect 4009 16294 4021 16346
rect 4021 16294 4051 16346
rect 4075 16294 4085 16346
rect 4085 16294 4131 16346
rect 3835 16292 3891 16294
rect 3915 16292 3971 16294
rect 3995 16292 4051 16294
rect 4075 16292 4131 16294
rect 3146 15308 3148 15328
rect 3148 15308 3200 15328
rect 3200 15308 3202 15328
rect 3146 15272 3202 15308
rect 4066 16088 4122 16144
rect 3175 14714 3231 14716
rect 3255 14714 3311 14716
rect 3335 14714 3391 14716
rect 3415 14714 3471 14716
rect 3175 14662 3221 14714
rect 3221 14662 3231 14714
rect 3255 14662 3285 14714
rect 3285 14662 3297 14714
rect 3297 14662 3311 14714
rect 3335 14662 3349 14714
rect 3349 14662 3361 14714
rect 3361 14662 3391 14714
rect 3415 14662 3425 14714
rect 3425 14662 3471 14714
rect 3175 14660 3231 14662
rect 3255 14660 3311 14662
rect 3335 14660 3391 14662
rect 3415 14660 3471 14662
rect 3835 15258 3891 15260
rect 3915 15258 3971 15260
rect 3995 15258 4051 15260
rect 4075 15258 4131 15260
rect 3835 15206 3881 15258
rect 3881 15206 3891 15258
rect 3915 15206 3945 15258
rect 3945 15206 3957 15258
rect 3957 15206 3971 15258
rect 3995 15206 4009 15258
rect 4009 15206 4021 15258
rect 4021 15206 4051 15258
rect 4075 15206 4085 15258
rect 4085 15206 4131 15258
rect 3835 15204 3891 15206
rect 3915 15204 3971 15206
rect 3995 15204 4051 15206
rect 4075 15204 4131 15206
rect 5262 16516 5318 16552
rect 5262 16496 5264 16516
rect 5264 16496 5316 16516
rect 5316 16496 5318 16516
rect 4618 15136 4674 15192
rect 4434 14900 4436 14920
rect 4436 14900 4488 14920
rect 4488 14900 4490 14920
rect 4434 14864 4490 14900
rect 3835 14170 3891 14172
rect 3915 14170 3971 14172
rect 3995 14170 4051 14172
rect 4075 14170 4131 14172
rect 3835 14118 3881 14170
rect 3881 14118 3891 14170
rect 3915 14118 3945 14170
rect 3945 14118 3957 14170
rect 3957 14118 3971 14170
rect 3995 14118 4009 14170
rect 4009 14118 4021 14170
rect 4021 14118 4051 14170
rect 4075 14118 4085 14170
rect 4085 14118 4131 14170
rect 3835 14116 3891 14118
rect 3915 14116 3971 14118
rect 3995 14116 4051 14118
rect 4075 14116 4131 14118
rect 3175 13626 3231 13628
rect 3255 13626 3311 13628
rect 3335 13626 3391 13628
rect 3415 13626 3471 13628
rect 3175 13574 3221 13626
rect 3221 13574 3231 13626
rect 3255 13574 3285 13626
rect 3285 13574 3297 13626
rect 3297 13574 3311 13626
rect 3335 13574 3349 13626
rect 3349 13574 3361 13626
rect 3361 13574 3391 13626
rect 3415 13574 3425 13626
rect 3425 13574 3471 13626
rect 3175 13572 3231 13574
rect 3255 13572 3311 13574
rect 3335 13572 3391 13574
rect 3415 13572 3471 13574
rect 2594 8336 2650 8392
rect 2410 6840 2466 6896
rect 2318 6160 2374 6216
rect 2686 7928 2742 7984
rect 2594 6160 2650 6216
rect 2594 5072 2650 5128
rect 3974 13504 4030 13560
rect 3606 13252 3662 13288
rect 3606 13232 3608 13252
rect 3608 13232 3660 13252
rect 3660 13232 3662 13252
rect 3835 13082 3891 13084
rect 3915 13082 3971 13084
rect 3995 13082 4051 13084
rect 4075 13082 4131 13084
rect 3835 13030 3881 13082
rect 3881 13030 3891 13082
rect 3915 13030 3945 13082
rect 3945 13030 3957 13082
rect 3957 13030 3971 13082
rect 3995 13030 4009 13082
rect 4009 13030 4021 13082
rect 4021 13030 4051 13082
rect 4075 13030 4085 13082
rect 4085 13030 4131 13082
rect 3835 13028 3891 13030
rect 3915 13028 3971 13030
rect 3995 13028 4051 13030
rect 4075 13028 4131 13030
rect 3175 12538 3231 12540
rect 3255 12538 3311 12540
rect 3335 12538 3391 12540
rect 3415 12538 3471 12540
rect 3175 12486 3221 12538
rect 3221 12486 3231 12538
rect 3255 12486 3285 12538
rect 3285 12486 3297 12538
rect 3297 12486 3311 12538
rect 3335 12486 3349 12538
rect 3349 12486 3361 12538
rect 3361 12486 3391 12538
rect 3415 12486 3425 12538
rect 3425 12486 3471 12538
rect 3175 12484 3231 12486
rect 3255 12484 3311 12486
rect 3335 12484 3391 12486
rect 3415 12484 3471 12486
rect 3175 11450 3231 11452
rect 3255 11450 3311 11452
rect 3335 11450 3391 11452
rect 3415 11450 3471 11452
rect 3175 11398 3221 11450
rect 3221 11398 3231 11450
rect 3255 11398 3285 11450
rect 3285 11398 3297 11450
rect 3297 11398 3311 11450
rect 3335 11398 3349 11450
rect 3349 11398 3361 11450
rect 3361 11398 3391 11450
rect 3415 11398 3425 11450
rect 3425 11398 3471 11450
rect 3175 11396 3231 11398
rect 3255 11396 3311 11398
rect 3335 11396 3391 11398
rect 3415 11396 3471 11398
rect 3330 10648 3386 10704
rect 3698 12416 3754 12472
rect 4342 14048 4398 14104
rect 4250 12960 4306 13016
rect 3835 11994 3891 11996
rect 3915 11994 3971 11996
rect 3995 11994 4051 11996
rect 4075 11994 4131 11996
rect 3835 11942 3881 11994
rect 3881 11942 3891 11994
rect 3915 11942 3945 11994
rect 3945 11942 3957 11994
rect 3957 11942 3971 11994
rect 3995 11942 4009 11994
rect 4009 11942 4021 11994
rect 4021 11942 4051 11994
rect 4075 11942 4085 11994
rect 4085 11942 4131 11994
rect 3835 11940 3891 11942
rect 3915 11940 3971 11942
rect 3995 11940 4051 11942
rect 4075 11940 4131 11942
rect 4250 12280 4306 12336
rect 3835 10906 3891 10908
rect 3915 10906 3971 10908
rect 3995 10906 4051 10908
rect 4075 10906 4131 10908
rect 3835 10854 3881 10906
rect 3881 10854 3891 10906
rect 3915 10854 3945 10906
rect 3945 10854 3957 10906
rect 3957 10854 3971 10906
rect 3995 10854 4009 10906
rect 4009 10854 4021 10906
rect 4021 10854 4051 10906
rect 4075 10854 4085 10906
rect 4085 10854 4131 10906
rect 3835 10852 3891 10854
rect 3915 10852 3971 10854
rect 3995 10852 4051 10854
rect 4075 10852 4131 10854
rect 3175 10362 3231 10364
rect 3255 10362 3311 10364
rect 3335 10362 3391 10364
rect 3415 10362 3471 10364
rect 3175 10310 3221 10362
rect 3221 10310 3231 10362
rect 3255 10310 3285 10362
rect 3285 10310 3297 10362
rect 3297 10310 3311 10362
rect 3335 10310 3349 10362
rect 3349 10310 3361 10362
rect 3361 10310 3391 10362
rect 3415 10310 3425 10362
rect 3425 10310 3471 10362
rect 3175 10308 3231 10310
rect 3255 10308 3311 10310
rect 3335 10308 3391 10310
rect 3415 10308 3471 10310
rect 3422 9580 3478 9616
rect 3422 9560 3424 9580
rect 3424 9560 3476 9580
rect 3476 9560 3478 9580
rect 3175 9274 3231 9276
rect 3255 9274 3311 9276
rect 3335 9274 3391 9276
rect 3415 9274 3471 9276
rect 3175 9222 3221 9274
rect 3221 9222 3231 9274
rect 3255 9222 3285 9274
rect 3285 9222 3297 9274
rect 3297 9222 3311 9274
rect 3335 9222 3349 9274
rect 3349 9222 3361 9274
rect 3361 9222 3391 9274
rect 3415 9222 3425 9274
rect 3425 9222 3471 9274
rect 3175 9220 3231 9222
rect 3255 9220 3311 9222
rect 3335 9220 3391 9222
rect 3415 9220 3471 9222
rect 2962 6296 3018 6352
rect 2962 4120 3018 4176
rect 3175 8186 3231 8188
rect 3255 8186 3311 8188
rect 3335 8186 3391 8188
rect 3415 8186 3471 8188
rect 3175 8134 3221 8186
rect 3221 8134 3231 8186
rect 3255 8134 3285 8186
rect 3285 8134 3297 8186
rect 3297 8134 3311 8186
rect 3335 8134 3349 8186
rect 3349 8134 3361 8186
rect 3361 8134 3391 8186
rect 3415 8134 3425 8186
rect 3425 8134 3471 8186
rect 3175 8132 3231 8134
rect 3255 8132 3311 8134
rect 3335 8132 3391 8134
rect 3415 8132 3471 8134
rect 3422 7928 3478 7984
rect 4066 10376 4122 10432
rect 3835 9818 3891 9820
rect 3915 9818 3971 9820
rect 3995 9818 4051 9820
rect 4075 9818 4131 9820
rect 3835 9766 3881 9818
rect 3881 9766 3891 9818
rect 3915 9766 3945 9818
rect 3945 9766 3957 9818
rect 3957 9766 3971 9818
rect 3995 9766 4009 9818
rect 4009 9766 4021 9818
rect 4021 9766 4051 9818
rect 4075 9766 4085 9818
rect 4085 9766 4131 9818
rect 3835 9764 3891 9766
rect 3915 9764 3971 9766
rect 3995 9764 4051 9766
rect 4075 9764 4131 9766
rect 4158 9560 4214 9616
rect 4250 9152 4306 9208
rect 4434 11736 4490 11792
rect 4250 8880 4306 8936
rect 3835 8730 3891 8732
rect 3915 8730 3971 8732
rect 3995 8730 4051 8732
rect 4075 8730 4131 8732
rect 3835 8678 3881 8730
rect 3881 8678 3891 8730
rect 3915 8678 3945 8730
rect 3945 8678 3957 8730
rect 3957 8678 3971 8730
rect 3995 8678 4009 8730
rect 4009 8678 4021 8730
rect 4021 8678 4051 8730
rect 4075 8678 4085 8730
rect 4085 8678 4131 8730
rect 3835 8676 3891 8678
rect 3915 8676 3971 8678
rect 3995 8676 4051 8678
rect 4075 8676 4131 8678
rect 3835 7642 3891 7644
rect 3915 7642 3971 7644
rect 3995 7642 4051 7644
rect 4075 7642 4131 7644
rect 3835 7590 3881 7642
rect 3881 7590 3891 7642
rect 3915 7590 3945 7642
rect 3945 7590 3957 7642
rect 3957 7590 3971 7642
rect 3995 7590 4009 7642
rect 4009 7590 4021 7642
rect 4021 7590 4051 7642
rect 4075 7590 4085 7642
rect 4085 7590 4131 7642
rect 3835 7588 3891 7590
rect 3915 7588 3971 7590
rect 3995 7588 4051 7590
rect 4075 7588 4131 7590
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 3422 6160 3478 6216
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 4066 6724 4122 6760
rect 4066 6704 4068 6724
rect 4068 6704 4120 6724
rect 4120 6704 4122 6724
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 3835 6554 3891 6556
rect 3915 6554 3971 6556
rect 3995 6554 4051 6556
rect 4075 6554 4131 6556
rect 3835 6502 3881 6554
rect 3881 6502 3891 6554
rect 3915 6502 3945 6554
rect 3945 6502 3957 6554
rect 3957 6502 3971 6554
rect 3995 6502 4009 6554
rect 4009 6502 4021 6554
rect 4021 6502 4051 6554
rect 4075 6502 4085 6554
rect 4085 6502 4131 6554
rect 3835 6500 3891 6502
rect 3915 6500 3971 6502
rect 3995 6500 4051 6502
rect 4075 6500 4131 6502
rect 4710 14184 4766 14240
rect 4618 11600 4674 11656
rect 4526 10784 4582 10840
rect 4710 11056 4766 11112
rect 4894 13812 4896 13832
rect 4896 13812 4948 13832
rect 4948 13812 4950 13832
rect 4894 13776 4950 13812
rect 4894 12144 4950 12200
rect 4526 8200 4582 8256
rect 4342 6976 4398 7032
rect 4710 8064 4766 8120
rect 4618 7248 4674 7304
rect 3835 5466 3891 5468
rect 3915 5466 3971 5468
rect 3995 5466 4051 5468
rect 4075 5466 4131 5468
rect 3835 5414 3881 5466
rect 3881 5414 3891 5466
rect 3915 5414 3945 5466
rect 3945 5414 3957 5466
rect 3957 5414 3971 5466
rect 3995 5414 4009 5466
rect 4009 5414 4021 5466
rect 4021 5414 4051 5466
rect 4075 5414 4085 5466
rect 4085 5414 4131 5466
rect 3835 5412 3891 5414
rect 3915 5412 3971 5414
rect 3995 5412 4051 5414
rect 4075 5412 4131 5414
rect 3882 5208 3938 5264
rect 4158 5208 4214 5264
rect 3835 4378 3891 4380
rect 3915 4378 3971 4380
rect 3995 4378 4051 4380
rect 4075 4378 4131 4380
rect 3835 4326 3881 4378
rect 3881 4326 3891 4378
rect 3915 4326 3945 4378
rect 3945 4326 3957 4378
rect 3957 4326 3971 4378
rect 3995 4326 4009 4378
rect 4009 4326 4021 4378
rect 4021 4326 4051 4378
rect 4075 4326 4085 4378
rect 4085 4326 4131 4378
rect 3835 4324 3891 4326
rect 3915 4324 3971 4326
rect 3995 4324 4051 4326
rect 4075 4324 4131 4326
rect 4434 4020 4436 4040
rect 4436 4020 4488 4040
rect 4488 4020 4490 4040
rect 4434 3984 4490 4020
rect 4434 3440 4490 3496
rect 5078 13132 5080 13152
rect 5080 13132 5132 13152
rect 5132 13132 5134 13152
rect 5078 13096 5134 13132
rect 5354 15020 5410 15056
rect 5354 15000 5356 15020
rect 5356 15000 5408 15020
rect 5408 15000 5410 15020
rect 5262 13504 5318 13560
rect 5170 12552 5226 12608
rect 5446 13640 5502 13696
rect 5446 13504 5502 13560
rect 5814 16632 5870 16688
rect 5998 15544 6054 15600
rect 5906 15408 5962 15464
rect 5906 15000 5962 15056
rect 5446 12008 5502 12064
rect 5170 11328 5226 11384
rect 5170 10784 5226 10840
rect 5170 7792 5226 7848
rect 5078 6840 5134 6896
rect 5170 6704 5226 6760
rect 3835 3290 3891 3292
rect 3915 3290 3971 3292
rect 3995 3290 4051 3292
rect 4075 3290 4131 3292
rect 3835 3238 3881 3290
rect 3881 3238 3891 3290
rect 3915 3238 3945 3290
rect 3945 3238 3957 3290
rect 3957 3238 3971 3290
rect 3995 3238 4009 3290
rect 4009 3238 4021 3290
rect 4021 3238 4051 3290
rect 4075 3238 4085 3290
rect 4085 3238 4131 3290
rect 3835 3236 3891 3238
rect 3915 3236 3971 3238
rect 3995 3236 4051 3238
rect 4075 3236 4131 3238
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 4986 4564 4988 4584
rect 4988 4564 5040 4584
rect 5040 4564 5042 4584
rect 4986 4528 5042 4564
rect 5170 4528 5226 4584
rect 5538 10784 5594 10840
rect 5446 9868 5448 9888
rect 5448 9868 5500 9888
rect 5500 9868 5502 9888
rect 5446 9832 5502 9868
rect 2134 2080 2190 2136
rect 846 1536 902 1592
rect 2778 720 2834 776
rect 5814 10920 5870 10976
rect 5630 7928 5686 7984
rect 5630 6432 5686 6488
rect 6274 13776 6330 13832
rect 6182 13504 6238 13560
rect 6090 12588 6092 12608
rect 6092 12588 6144 12608
rect 6144 12588 6146 12608
rect 6090 12552 6146 12588
rect 15382 17992 15438 18048
rect 8022 17720 8078 17776
rect 6826 17332 6882 17368
rect 6826 17312 6828 17332
rect 6828 17312 6880 17332
rect 6880 17312 6882 17332
rect 7654 17312 7710 17368
rect 7286 17176 7342 17232
rect 6826 15816 6882 15872
rect 7614 16890 7670 16892
rect 7694 16890 7750 16892
rect 7774 16890 7830 16892
rect 7854 16890 7910 16892
rect 7614 16838 7660 16890
rect 7660 16838 7670 16890
rect 7694 16838 7724 16890
rect 7724 16838 7736 16890
rect 7736 16838 7750 16890
rect 7774 16838 7788 16890
rect 7788 16838 7800 16890
rect 7800 16838 7830 16890
rect 7854 16838 7864 16890
rect 7864 16838 7910 16890
rect 7614 16836 7670 16838
rect 7694 16836 7750 16838
rect 7774 16836 7830 16838
rect 7854 16836 7910 16838
rect 7286 16496 7342 16552
rect 7194 16224 7250 16280
rect 7614 15802 7670 15804
rect 7694 15802 7750 15804
rect 7774 15802 7830 15804
rect 7854 15802 7910 15804
rect 7614 15750 7660 15802
rect 7660 15750 7670 15802
rect 7694 15750 7724 15802
rect 7724 15750 7736 15802
rect 7736 15750 7750 15802
rect 7774 15750 7788 15802
rect 7788 15750 7800 15802
rect 7800 15750 7830 15802
rect 7854 15750 7864 15802
rect 7864 15750 7910 15802
rect 7614 15748 7670 15750
rect 7694 15748 7750 15750
rect 7774 15748 7830 15750
rect 7854 15748 7910 15750
rect 8274 17434 8330 17436
rect 8354 17434 8410 17436
rect 8434 17434 8490 17436
rect 8514 17434 8570 17436
rect 8274 17382 8320 17434
rect 8320 17382 8330 17434
rect 8354 17382 8384 17434
rect 8384 17382 8396 17434
rect 8396 17382 8410 17434
rect 8434 17382 8448 17434
rect 8448 17382 8460 17434
rect 8460 17382 8490 17434
rect 8514 17382 8524 17434
rect 8524 17382 8570 17434
rect 8274 17380 8330 17382
rect 8354 17380 8410 17382
rect 8434 17380 8490 17382
rect 8514 17380 8570 17382
rect 12713 17434 12769 17436
rect 12793 17434 12849 17436
rect 12873 17434 12929 17436
rect 12953 17434 13009 17436
rect 12713 17382 12759 17434
rect 12759 17382 12769 17434
rect 12793 17382 12823 17434
rect 12823 17382 12835 17434
rect 12835 17382 12849 17434
rect 12873 17382 12887 17434
rect 12887 17382 12899 17434
rect 12899 17382 12929 17434
rect 12953 17382 12963 17434
rect 12963 17382 13009 17434
rect 12713 17380 12769 17382
rect 12793 17380 12849 17382
rect 12873 17380 12929 17382
rect 12953 17380 13009 17382
rect 8390 16632 8446 16688
rect 8274 16346 8330 16348
rect 8354 16346 8410 16348
rect 8434 16346 8490 16348
rect 8514 16346 8570 16348
rect 8274 16294 8320 16346
rect 8320 16294 8330 16346
rect 8354 16294 8384 16346
rect 8384 16294 8396 16346
rect 8396 16294 8410 16346
rect 8434 16294 8448 16346
rect 8448 16294 8460 16346
rect 8460 16294 8490 16346
rect 8514 16294 8524 16346
rect 8524 16294 8570 16346
rect 8274 16292 8330 16294
rect 8354 16292 8410 16294
rect 8434 16292 8490 16294
rect 8514 16292 8570 16294
rect 8482 15972 8538 16008
rect 8482 15952 8484 15972
rect 8484 15952 8536 15972
rect 8536 15952 8538 15972
rect 8206 15852 8208 15872
rect 8208 15852 8260 15872
rect 8260 15852 8262 15872
rect 8206 15816 8262 15852
rect 8274 15258 8330 15260
rect 8354 15258 8410 15260
rect 8434 15258 8490 15260
rect 8514 15258 8570 15260
rect 8274 15206 8320 15258
rect 8320 15206 8330 15258
rect 8354 15206 8384 15258
rect 8384 15206 8396 15258
rect 8396 15206 8410 15258
rect 8434 15206 8448 15258
rect 8448 15206 8460 15258
rect 8460 15206 8490 15258
rect 8514 15206 8524 15258
rect 8524 15206 8570 15258
rect 8274 15204 8330 15206
rect 8354 15204 8410 15206
rect 8434 15204 8490 15206
rect 8514 15204 8570 15206
rect 8850 15816 8906 15872
rect 7102 14048 7158 14104
rect 6918 13640 6974 13696
rect 6182 9424 6238 9480
rect 5538 5480 5594 5536
rect 6458 10376 6514 10432
rect 6274 6840 6330 6896
rect 6826 12008 6882 12064
rect 6734 10920 6790 10976
rect 6642 10648 6698 10704
rect 6642 10104 6698 10160
rect 6918 9968 6974 10024
rect 6918 9424 6974 9480
rect 7286 11076 7342 11112
rect 7286 11056 7288 11076
rect 7288 11056 7340 11076
rect 7340 11056 7342 11076
rect 7930 14864 7986 14920
rect 7614 14714 7670 14716
rect 7694 14714 7750 14716
rect 7774 14714 7830 14716
rect 7854 14714 7910 14716
rect 7614 14662 7660 14714
rect 7660 14662 7670 14714
rect 7694 14662 7724 14714
rect 7724 14662 7736 14714
rect 7736 14662 7750 14714
rect 7774 14662 7788 14714
rect 7788 14662 7800 14714
rect 7800 14662 7830 14714
rect 7854 14662 7864 14714
rect 7864 14662 7910 14714
rect 7614 14660 7670 14662
rect 7694 14660 7750 14662
rect 7774 14660 7830 14662
rect 7854 14660 7910 14662
rect 8206 14592 8262 14648
rect 8114 14456 8170 14512
rect 8482 14456 8538 14512
rect 9126 16224 9182 16280
rect 9402 16904 9458 16960
rect 9126 15952 9182 16008
rect 9126 15272 9182 15328
rect 9034 14864 9090 14920
rect 8114 14184 8170 14240
rect 8022 13640 8078 13696
rect 7614 13626 7670 13628
rect 7694 13626 7750 13628
rect 7774 13626 7830 13628
rect 7854 13626 7910 13628
rect 7614 13574 7660 13626
rect 7660 13574 7670 13626
rect 7694 13574 7724 13626
rect 7724 13574 7736 13626
rect 7736 13574 7750 13626
rect 7774 13574 7788 13626
rect 7788 13574 7800 13626
rect 7800 13574 7830 13626
rect 7854 13574 7864 13626
rect 7864 13574 7910 13626
rect 7614 13572 7670 13574
rect 7694 13572 7750 13574
rect 7774 13572 7830 13574
rect 7854 13572 7910 13574
rect 8274 14170 8330 14172
rect 8354 14170 8410 14172
rect 8434 14170 8490 14172
rect 8514 14170 8570 14172
rect 8274 14118 8320 14170
rect 8320 14118 8330 14170
rect 8354 14118 8384 14170
rect 8384 14118 8396 14170
rect 8396 14118 8410 14170
rect 8434 14118 8448 14170
rect 8448 14118 8460 14170
rect 8460 14118 8490 14170
rect 8514 14118 8524 14170
rect 8524 14118 8570 14170
rect 8274 14116 8330 14118
rect 8354 14116 8410 14118
rect 8434 14116 8490 14118
rect 8514 14116 8570 14118
rect 8758 13912 8814 13968
rect 7562 12960 7618 13016
rect 8274 13082 8330 13084
rect 8354 13082 8410 13084
rect 8434 13082 8490 13084
rect 8514 13082 8570 13084
rect 8274 13030 8320 13082
rect 8320 13030 8330 13082
rect 8354 13030 8384 13082
rect 8384 13030 8396 13082
rect 8396 13030 8410 13082
rect 8434 13030 8448 13082
rect 8448 13030 8460 13082
rect 8460 13030 8490 13082
rect 8514 13030 8524 13082
rect 8524 13030 8570 13082
rect 8274 13028 8330 13030
rect 8354 13028 8410 13030
rect 8434 13028 8490 13030
rect 8514 13028 8570 13030
rect 7614 12538 7670 12540
rect 7694 12538 7750 12540
rect 7774 12538 7830 12540
rect 7854 12538 7910 12540
rect 7614 12486 7660 12538
rect 7660 12486 7670 12538
rect 7694 12486 7724 12538
rect 7724 12486 7736 12538
rect 7736 12486 7750 12538
rect 7774 12486 7788 12538
rect 7788 12486 7800 12538
rect 7800 12486 7830 12538
rect 7854 12486 7864 12538
rect 7864 12486 7910 12538
rect 7614 12484 7670 12486
rect 7694 12484 7750 12486
rect 7774 12484 7830 12486
rect 7854 12484 7910 12486
rect 8482 12688 8538 12744
rect 7746 11872 7802 11928
rect 8114 12280 8170 12336
rect 8022 12008 8078 12064
rect 7614 11450 7670 11452
rect 7694 11450 7750 11452
rect 7774 11450 7830 11452
rect 7854 11450 7910 11452
rect 7614 11398 7660 11450
rect 7660 11398 7670 11450
rect 7694 11398 7724 11450
rect 7724 11398 7736 11450
rect 7736 11398 7750 11450
rect 7774 11398 7788 11450
rect 7788 11398 7800 11450
rect 7800 11398 7830 11450
rect 7854 11398 7864 11450
rect 7864 11398 7910 11450
rect 7614 11396 7670 11398
rect 7694 11396 7750 11398
rect 7774 11396 7830 11398
rect 7854 11396 7910 11398
rect 7654 10920 7710 10976
rect 7746 10804 7802 10840
rect 7746 10784 7748 10804
rect 7748 10784 7800 10804
rect 7800 10784 7802 10804
rect 7378 10240 7434 10296
rect 7614 10362 7670 10364
rect 7694 10362 7750 10364
rect 7774 10362 7830 10364
rect 7854 10362 7910 10364
rect 7614 10310 7660 10362
rect 7660 10310 7670 10362
rect 7694 10310 7724 10362
rect 7724 10310 7736 10362
rect 7736 10310 7750 10362
rect 7774 10310 7788 10362
rect 7788 10310 7800 10362
rect 7800 10310 7830 10362
rect 7854 10310 7864 10362
rect 7864 10310 7910 10362
rect 7614 10308 7670 10310
rect 7694 10308 7750 10310
rect 7774 10308 7830 10310
rect 7854 10308 7910 10310
rect 7194 9832 7250 9888
rect 7654 9968 7710 10024
rect 7614 9274 7670 9276
rect 7694 9274 7750 9276
rect 7774 9274 7830 9276
rect 7854 9274 7910 9276
rect 7614 9222 7660 9274
rect 7660 9222 7670 9274
rect 7694 9222 7724 9274
rect 7724 9222 7736 9274
rect 7736 9222 7750 9274
rect 7774 9222 7788 9274
rect 7788 9222 7800 9274
rect 7800 9222 7830 9274
rect 7854 9222 7864 9274
rect 7864 9222 7910 9274
rect 7614 9220 7670 9222
rect 7694 9220 7750 9222
rect 7774 9220 7830 9222
rect 7854 9220 7910 9222
rect 6918 8472 6974 8528
rect 6918 8336 6974 8392
rect 7286 8608 7342 8664
rect 7102 8084 7158 8120
rect 7102 8064 7104 8084
rect 7104 8064 7156 8084
rect 7156 8064 7158 8084
rect 7102 7928 7158 7984
rect 7010 6568 7066 6624
rect 7010 6432 7066 6488
rect 6274 5616 6330 5672
rect 6090 5208 6146 5264
rect 5630 3476 5632 3496
rect 5632 3476 5684 3496
rect 5684 3476 5686 3496
rect 5630 3440 5686 3476
rect 6090 3460 6146 3496
rect 6090 3440 6092 3460
rect 6092 3440 6144 3460
rect 6144 3440 6146 3460
rect 6458 3732 6514 3768
rect 6458 3712 6460 3732
rect 6460 3712 6512 3732
rect 6512 3712 6514 3732
rect 6918 6024 6974 6080
rect 7838 8744 7894 8800
rect 7746 8336 7802 8392
rect 7614 8186 7670 8188
rect 7694 8186 7750 8188
rect 7774 8186 7830 8188
rect 7854 8186 7910 8188
rect 7614 8134 7660 8186
rect 7660 8134 7670 8186
rect 7694 8134 7724 8186
rect 7724 8134 7736 8186
rect 7736 8134 7750 8186
rect 7774 8134 7788 8186
rect 7788 8134 7800 8186
rect 7800 8134 7830 8186
rect 7854 8134 7864 8186
rect 7864 8134 7910 8186
rect 7614 8132 7670 8134
rect 7694 8132 7750 8134
rect 7774 8132 7830 8134
rect 7854 8132 7910 8134
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 7470 6840 7526 6896
rect 7654 6568 7710 6624
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 7470 5208 7526 5264
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 7838 3576 7894 3632
rect 8274 11994 8330 11996
rect 8354 11994 8410 11996
rect 8434 11994 8490 11996
rect 8514 11994 8570 11996
rect 8274 11942 8320 11994
rect 8320 11942 8330 11994
rect 8354 11942 8384 11994
rect 8384 11942 8396 11994
rect 8396 11942 8410 11994
rect 8434 11942 8448 11994
rect 8448 11942 8460 11994
rect 8460 11942 8490 11994
rect 8514 11942 8524 11994
rect 8524 11942 8570 11994
rect 8274 11940 8330 11942
rect 8354 11940 8410 11942
rect 8434 11940 8490 11942
rect 8514 11940 8570 11942
rect 8390 11328 8446 11384
rect 8274 10906 8330 10908
rect 8354 10906 8410 10908
rect 8434 10906 8490 10908
rect 8514 10906 8570 10908
rect 8274 10854 8320 10906
rect 8320 10854 8330 10906
rect 8354 10854 8384 10906
rect 8384 10854 8396 10906
rect 8396 10854 8410 10906
rect 8434 10854 8448 10906
rect 8448 10854 8460 10906
rect 8460 10854 8490 10906
rect 8514 10854 8524 10906
rect 8524 10854 8570 10906
rect 8274 10852 8330 10854
rect 8354 10852 8410 10854
rect 8434 10852 8490 10854
rect 8514 10852 8570 10854
rect 8574 10668 8630 10704
rect 8574 10648 8576 10668
rect 8576 10648 8628 10668
rect 8628 10648 8630 10668
rect 8482 10376 8538 10432
rect 8298 10104 8354 10160
rect 8206 10004 8208 10024
rect 8208 10004 8260 10024
rect 8260 10004 8262 10024
rect 8206 9968 8262 10004
rect 8274 9818 8330 9820
rect 8354 9818 8410 9820
rect 8434 9818 8490 9820
rect 8514 9818 8570 9820
rect 8274 9766 8320 9818
rect 8320 9766 8330 9818
rect 8354 9766 8384 9818
rect 8384 9766 8396 9818
rect 8396 9766 8410 9818
rect 8434 9766 8448 9818
rect 8448 9766 8460 9818
rect 8460 9766 8490 9818
rect 8514 9766 8524 9818
rect 8524 9766 8570 9818
rect 8274 9764 8330 9766
rect 8354 9764 8410 9766
rect 8434 9764 8490 9766
rect 8514 9764 8570 9766
rect 8758 12960 8814 13016
rect 8942 13776 8998 13832
rect 8390 9152 8446 9208
rect 8850 9832 8906 9888
rect 8274 8730 8330 8732
rect 8354 8730 8410 8732
rect 8434 8730 8490 8732
rect 8514 8730 8570 8732
rect 8274 8678 8320 8730
rect 8320 8678 8330 8730
rect 8354 8678 8384 8730
rect 8384 8678 8396 8730
rect 8396 8678 8410 8730
rect 8434 8678 8448 8730
rect 8448 8678 8460 8730
rect 8460 8678 8490 8730
rect 8514 8678 8524 8730
rect 8524 8678 8570 8730
rect 8274 8676 8330 8678
rect 8354 8676 8410 8678
rect 8434 8676 8490 8678
rect 8514 8676 8570 8678
rect 8114 8608 8170 8664
rect 8114 8336 8170 8392
rect 8274 7642 8330 7644
rect 8354 7642 8410 7644
rect 8434 7642 8490 7644
rect 8514 7642 8570 7644
rect 8274 7590 8320 7642
rect 8320 7590 8330 7642
rect 8354 7590 8384 7642
rect 8384 7590 8396 7642
rect 8396 7590 8410 7642
rect 8434 7590 8448 7642
rect 8448 7590 8460 7642
rect 8460 7590 8490 7642
rect 8514 7590 8524 7642
rect 8524 7590 8570 7642
rect 8274 7588 8330 7590
rect 8354 7588 8410 7590
rect 8434 7588 8490 7590
rect 8514 7588 8570 7590
rect 8274 6554 8330 6556
rect 8354 6554 8410 6556
rect 8434 6554 8490 6556
rect 8514 6554 8570 6556
rect 8274 6502 8320 6554
rect 8320 6502 8330 6554
rect 8354 6502 8384 6554
rect 8384 6502 8396 6554
rect 8396 6502 8410 6554
rect 8434 6502 8448 6554
rect 8448 6502 8460 6554
rect 8460 6502 8490 6554
rect 8514 6502 8524 6554
rect 8524 6502 8570 6554
rect 8274 6500 8330 6502
rect 8354 6500 8410 6502
rect 8434 6500 8490 6502
rect 8514 6500 8570 6502
rect 8022 5888 8078 5944
rect 8022 5108 8024 5128
rect 8024 5108 8076 5128
rect 8076 5108 8078 5128
rect 8022 5072 8078 5108
rect 8022 4800 8078 4856
rect 8022 4392 8078 4448
rect 8022 3984 8078 4040
rect 8482 5888 8538 5944
rect 8206 5616 8262 5672
rect 8666 5888 8722 5944
rect 8274 5466 8330 5468
rect 8354 5466 8410 5468
rect 8434 5466 8490 5468
rect 8514 5466 8570 5468
rect 8274 5414 8320 5466
rect 8320 5414 8330 5466
rect 8354 5414 8384 5466
rect 8384 5414 8396 5466
rect 8396 5414 8410 5466
rect 8434 5414 8448 5466
rect 8448 5414 8460 5466
rect 8460 5414 8490 5466
rect 8514 5414 8524 5466
rect 8524 5414 8570 5466
rect 8274 5412 8330 5414
rect 8354 5412 8410 5414
rect 8434 5412 8490 5414
rect 8514 5412 8570 5414
rect 8274 4378 8330 4380
rect 8354 4378 8410 4380
rect 8434 4378 8490 4380
rect 8514 4378 8570 4380
rect 8274 4326 8320 4378
rect 8320 4326 8330 4378
rect 8354 4326 8384 4378
rect 8384 4326 8396 4378
rect 8396 4326 8410 4378
rect 8434 4326 8448 4378
rect 8448 4326 8460 4378
rect 8460 4326 8490 4378
rect 8514 4326 8524 4378
rect 8524 4326 8570 4378
rect 8274 4324 8330 4326
rect 8354 4324 8410 4326
rect 8434 4324 8490 4326
rect 8514 4324 8570 4326
rect 9402 15408 9458 15464
rect 9586 16224 9642 16280
rect 9586 15408 9642 15464
rect 9494 13912 9550 13968
rect 9218 13096 9274 13152
rect 9218 12552 9274 12608
rect 9034 10648 9090 10704
rect 9218 11892 9274 11928
rect 9218 11872 9220 11892
rect 9220 11872 9272 11892
rect 9272 11872 9274 11892
rect 10046 14456 10102 14512
rect 9678 12416 9734 12472
rect 9126 9560 9182 9616
rect 9586 11600 9642 11656
rect 9402 10648 9458 10704
rect 9310 10260 9366 10296
rect 9310 10240 9312 10260
rect 9312 10240 9364 10260
rect 9364 10240 9366 10260
rect 9126 8336 9182 8392
rect 9126 8200 9182 8256
rect 9034 7692 9036 7712
rect 9036 7692 9088 7712
rect 9088 7692 9090 7712
rect 9034 7656 9090 7692
rect 9034 7384 9090 7440
rect 9770 10240 9826 10296
rect 9586 9016 9642 9072
rect 9402 8064 9458 8120
rect 9494 6432 9550 6488
rect 9402 4664 9458 4720
rect 8274 3290 8330 3292
rect 8354 3290 8410 3292
rect 8434 3290 8490 3292
rect 8514 3290 8570 3292
rect 8274 3238 8320 3290
rect 8320 3238 8330 3290
rect 8354 3238 8384 3290
rect 8384 3238 8396 3290
rect 8396 3238 8410 3290
rect 8434 3238 8448 3290
rect 8448 3238 8460 3290
rect 8460 3238 8490 3290
rect 8514 3238 8524 3290
rect 8524 3238 8570 3290
rect 8274 3236 8330 3238
rect 8354 3236 8410 3238
rect 8434 3236 8490 3238
rect 8514 3236 8570 3238
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 3835 2202 3891 2204
rect 3915 2202 3971 2204
rect 3995 2202 4051 2204
rect 4075 2202 4131 2204
rect 3835 2150 3881 2202
rect 3881 2150 3891 2202
rect 3915 2150 3945 2202
rect 3945 2150 3957 2202
rect 3957 2150 3971 2202
rect 3995 2150 4009 2202
rect 4009 2150 4021 2202
rect 4021 2150 4051 2202
rect 4075 2150 4085 2202
rect 4085 2150 4131 2202
rect 3835 2148 3891 2150
rect 3915 2148 3971 2150
rect 3995 2148 4051 2150
rect 4075 2148 4131 2150
rect 10230 14456 10286 14512
rect 10138 13096 10194 13152
rect 10414 12552 10470 12608
rect 10414 12280 10470 12336
rect 10046 11600 10102 11656
rect 10046 10512 10102 10568
rect 9862 6568 9918 6624
rect 10322 11464 10378 11520
rect 10506 11328 10562 11384
rect 10230 10648 10286 10704
rect 10322 10240 10378 10296
rect 10230 9560 10286 9616
rect 10138 9152 10194 9208
rect 8274 2202 8330 2204
rect 8354 2202 8410 2204
rect 8434 2202 8490 2204
rect 8514 2202 8570 2204
rect 8274 2150 8320 2202
rect 8320 2150 8330 2202
rect 8354 2150 8384 2202
rect 8384 2150 8396 2202
rect 8396 2150 8410 2202
rect 8434 2150 8448 2202
rect 8448 2150 8460 2202
rect 8460 2150 8490 2202
rect 8514 2150 8524 2202
rect 8524 2150 8570 2202
rect 8274 2148 8330 2150
rect 8354 2148 8410 2150
rect 8434 2148 8490 2150
rect 8514 2148 8570 2150
rect 2870 40 2926 96
rect 10046 5208 10102 5264
rect 10322 5788 10324 5808
rect 10324 5788 10376 5808
rect 10376 5788 10378 5808
rect 10322 5752 10378 5788
rect 10322 4120 10378 4176
rect 10966 16632 11022 16688
rect 10782 14184 10838 14240
rect 10966 15136 11022 15192
rect 12346 17176 12402 17232
rect 12162 17040 12218 17096
rect 12053 16890 12109 16892
rect 12133 16890 12189 16892
rect 12213 16890 12269 16892
rect 12293 16890 12349 16892
rect 12053 16838 12099 16890
rect 12099 16838 12109 16890
rect 12133 16838 12163 16890
rect 12163 16838 12175 16890
rect 12175 16838 12189 16890
rect 12213 16838 12227 16890
rect 12227 16838 12239 16890
rect 12239 16838 12269 16890
rect 12293 16838 12303 16890
rect 12303 16838 12349 16890
rect 12053 16836 12109 16838
rect 12133 16836 12189 16838
rect 12213 16836 12269 16838
rect 12293 16836 12349 16838
rect 11242 16632 11298 16688
rect 11242 13252 11298 13288
rect 11242 13232 11244 13252
rect 11244 13232 11296 13252
rect 11296 13232 11298 13252
rect 10782 10140 10784 10160
rect 10784 10140 10836 10160
rect 10836 10140 10838 10160
rect 10782 10104 10838 10140
rect 11058 12180 11060 12200
rect 11060 12180 11112 12200
rect 11112 12180 11114 12200
rect 11058 12144 11114 12180
rect 10966 10376 11022 10432
rect 11058 8608 11114 8664
rect 11334 12552 11390 12608
rect 11334 11772 11336 11792
rect 11336 11772 11388 11792
rect 11388 11772 11390 11792
rect 11334 11736 11390 11772
rect 11242 10648 11298 10704
rect 11242 9596 11244 9616
rect 11244 9596 11296 9616
rect 11296 9596 11298 9616
rect 11242 9560 11298 9596
rect 11242 9152 11298 9208
rect 10598 5480 10654 5536
rect 10966 6160 11022 6216
rect 12530 16244 12586 16280
rect 12530 16224 12532 16244
rect 12532 16224 12584 16244
rect 12584 16224 12586 16244
rect 12053 15802 12109 15804
rect 12133 15802 12189 15804
rect 12213 15802 12269 15804
rect 12293 15802 12349 15804
rect 12053 15750 12099 15802
rect 12099 15750 12109 15802
rect 12133 15750 12163 15802
rect 12163 15750 12175 15802
rect 12175 15750 12189 15802
rect 12213 15750 12227 15802
rect 12227 15750 12239 15802
rect 12239 15750 12269 15802
rect 12293 15750 12303 15802
rect 12303 15750 12349 15802
rect 12053 15748 12109 15750
rect 12133 15748 12189 15750
rect 12213 15748 12269 15750
rect 12293 15748 12349 15750
rect 12530 15544 12586 15600
rect 12070 15272 12126 15328
rect 12438 15000 12494 15056
rect 12438 14728 12494 14784
rect 12053 14714 12109 14716
rect 12133 14714 12189 14716
rect 12213 14714 12269 14716
rect 12293 14714 12349 14716
rect 12053 14662 12099 14714
rect 12099 14662 12109 14714
rect 12133 14662 12163 14714
rect 12163 14662 12175 14714
rect 12175 14662 12189 14714
rect 12213 14662 12227 14714
rect 12227 14662 12239 14714
rect 12239 14662 12269 14714
rect 12293 14662 12303 14714
rect 12303 14662 12349 14714
rect 12053 14660 12109 14662
rect 12133 14660 12189 14662
rect 12213 14660 12269 14662
rect 12293 14660 12349 14662
rect 12713 16346 12769 16348
rect 12793 16346 12849 16348
rect 12873 16346 12929 16348
rect 12953 16346 13009 16348
rect 12713 16294 12759 16346
rect 12759 16294 12769 16346
rect 12793 16294 12823 16346
rect 12823 16294 12835 16346
rect 12835 16294 12849 16346
rect 12873 16294 12887 16346
rect 12887 16294 12899 16346
rect 12899 16294 12929 16346
rect 12953 16294 12963 16346
rect 12963 16294 13009 16346
rect 12713 16292 12769 16294
rect 12793 16292 12849 16294
rect 12873 16292 12929 16294
rect 12953 16292 13009 16294
rect 12714 16108 12770 16144
rect 12714 16088 12716 16108
rect 12716 16088 12768 16108
rect 12768 16088 12770 16108
rect 12713 15258 12769 15260
rect 12793 15258 12849 15260
rect 12873 15258 12929 15260
rect 12953 15258 13009 15260
rect 12713 15206 12759 15258
rect 12759 15206 12769 15258
rect 12793 15206 12823 15258
rect 12823 15206 12835 15258
rect 12835 15206 12849 15258
rect 12873 15206 12887 15258
rect 12887 15206 12899 15258
rect 12899 15206 12929 15258
rect 12953 15206 12963 15258
rect 12963 15206 13009 15258
rect 12713 15204 12769 15206
rect 12793 15204 12849 15206
rect 12873 15204 12929 15206
rect 12953 15204 13009 15206
rect 11794 13640 11850 13696
rect 12053 13626 12109 13628
rect 12133 13626 12189 13628
rect 12213 13626 12269 13628
rect 12293 13626 12349 13628
rect 12053 13574 12099 13626
rect 12099 13574 12109 13626
rect 12133 13574 12163 13626
rect 12163 13574 12175 13626
rect 12175 13574 12189 13626
rect 12213 13574 12227 13626
rect 12227 13574 12239 13626
rect 12239 13574 12269 13626
rect 12293 13574 12303 13626
rect 12303 13574 12349 13626
rect 12053 13572 12109 13574
rect 12133 13572 12189 13574
rect 12213 13572 12269 13574
rect 12293 13572 12349 13574
rect 12070 13268 12072 13288
rect 12072 13268 12124 13288
rect 12124 13268 12126 13288
rect 12070 13232 12126 13268
rect 11794 12824 11850 12880
rect 11702 10240 11758 10296
rect 11518 9696 11574 9752
rect 12254 12688 12310 12744
rect 12053 12538 12109 12540
rect 12133 12538 12189 12540
rect 12213 12538 12269 12540
rect 12293 12538 12349 12540
rect 12053 12486 12099 12538
rect 12099 12486 12109 12538
rect 12133 12486 12163 12538
rect 12163 12486 12175 12538
rect 12175 12486 12189 12538
rect 12213 12486 12227 12538
rect 12227 12486 12239 12538
rect 12239 12486 12269 12538
rect 12293 12486 12303 12538
rect 12303 12486 12349 12538
rect 12053 12484 12109 12486
rect 12133 12484 12189 12486
rect 12213 12484 12269 12486
rect 12293 12484 12349 12486
rect 12713 14170 12769 14172
rect 12793 14170 12849 14172
rect 12873 14170 12929 14172
rect 12953 14170 13009 14172
rect 12713 14118 12759 14170
rect 12759 14118 12769 14170
rect 12793 14118 12823 14170
rect 12823 14118 12835 14170
rect 12835 14118 12849 14170
rect 12873 14118 12887 14170
rect 12887 14118 12899 14170
rect 12899 14118 12929 14170
rect 12953 14118 12963 14170
rect 12963 14118 13009 14170
rect 12713 14116 12769 14118
rect 12793 14116 12849 14118
rect 12873 14116 12929 14118
rect 12953 14116 13009 14118
rect 12898 13912 12954 13968
rect 12713 13082 12769 13084
rect 12793 13082 12849 13084
rect 12873 13082 12929 13084
rect 12953 13082 13009 13084
rect 12713 13030 12759 13082
rect 12759 13030 12769 13082
rect 12793 13030 12823 13082
rect 12823 13030 12835 13082
rect 12835 13030 12849 13082
rect 12873 13030 12887 13082
rect 12887 13030 12899 13082
rect 12899 13030 12929 13082
rect 12953 13030 12963 13082
rect 12963 13030 13009 13082
rect 12713 13028 12769 13030
rect 12793 13028 12849 13030
rect 12873 13028 12929 13030
rect 12953 13028 13009 13030
rect 12806 12688 12862 12744
rect 13082 12416 13138 12472
rect 12438 12280 12494 12336
rect 12438 11872 12494 11928
rect 12438 11464 12494 11520
rect 12053 11450 12109 11452
rect 12133 11450 12189 11452
rect 12213 11450 12269 11452
rect 12293 11450 12349 11452
rect 12053 11398 12099 11450
rect 12099 11398 12109 11450
rect 12133 11398 12163 11450
rect 12163 11398 12175 11450
rect 12175 11398 12189 11450
rect 12213 11398 12227 11450
rect 12227 11398 12239 11450
rect 12239 11398 12269 11450
rect 12293 11398 12303 11450
rect 12303 11398 12349 11450
rect 12053 11396 12109 11398
rect 12133 11396 12189 11398
rect 12213 11396 12269 11398
rect 12293 11396 12349 11398
rect 12438 10784 12494 10840
rect 12438 10648 12494 10704
rect 12438 10376 12494 10432
rect 12053 10362 12109 10364
rect 12133 10362 12189 10364
rect 12213 10362 12269 10364
rect 12293 10362 12349 10364
rect 12053 10310 12099 10362
rect 12099 10310 12109 10362
rect 12133 10310 12163 10362
rect 12163 10310 12175 10362
rect 12175 10310 12189 10362
rect 12213 10310 12227 10362
rect 12227 10310 12239 10362
rect 12239 10310 12269 10362
rect 12293 10310 12303 10362
rect 12303 10310 12349 10362
rect 12053 10308 12109 10310
rect 12133 10308 12189 10310
rect 12213 10308 12269 10310
rect 12293 10308 12349 10310
rect 12438 10240 12494 10296
rect 11702 9560 11758 9616
rect 11886 9560 11942 9616
rect 11610 8780 11612 8800
rect 11612 8780 11664 8800
rect 11664 8780 11666 8800
rect 11610 8744 11666 8780
rect 11518 7520 11574 7576
rect 11794 9152 11850 9208
rect 10690 3052 10746 3088
rect 10690 3032 10692 3052
rect 10692 3032 10744 3052
rect 10744 3032 10746 3052
rect 11242 2896 11298 2952
rect 12713 11994 12769 11996
rect 12793 11994 12849 11996
rect 12873 11994 12929 11996
rect 12953 11994 13009 11996
rect 12713 11942 12759 11994
rect 12759 11942 12769 11994
rect 12793 11942 12823 11994
rect 12823 11942 12835 11994
rect 12835 11942 12849 11994
rect 12873 11942 12887 11994
rect 12887 11942 12899 11994
rect 12899 11942 12929 11994
rect 12953 11942 12963 11994
rect 12963 11942 13009 11994
rect 12713 11940 12769 11942
rect 12793 11940 12849 11942
rect 12873 11940 12929 11942
rect 12953 11940 13009 11942
rect 12898 11736 12954 11792
rect 12713 10906 12769 10908
rect 12793 10906 12849 10908
rect 12873 10906 12929 10908
rect 12953 10906 13009 10908
rect 12713 10854 12759 10906
rect 12759 10854 12769 10906
rect 12793 10854 12823 10906
rect 12823 10854 12835 10906
rect 12835 10854 12849 10906
rect 12873 10854 12887 10906
rect 12887 10854 12899 10906
rect 12899 10854 12929 10906
rect 12953 10854 12963 10906
rect 12963 10854 13009 10906
rect 12713 10852 12769 10854
rect 12793 10852 12849 10854
rect 12873 10852 12929 10854
rect 12953 10852 13009 10854
rect 12806 10104 12862 10160
rect 12990 10104 13046 10160
rect 14370 17584 14426 17640
rect 14278 15408 14334 15464
rect 14094 14864 14150 14920
rect 13726 13776 13782 13832
rect 13818 13368 13874 13424
rect 13910 13096 13966 13152
rect 14554 15272 14610 15328
rect 14186 13640 14242 13696
rect 14094 13096 14150 13152
rect 13450 11872 13506 11928
rect 13358 11464 13414 11520
rect 13358 11056 13414 11112
rect 13266 10784 13322 10840
rect 12713 9818 12769 9820
rect 12793 9818 12849 9820
rect 12873 9818 12929 9820
rect 12953 9818 13009 9820
rect 12713 9766 12759 9818
rect 12759 9766 12769 9818
rect 12793 9766 12823 9818
rect 12823 9766 12835 9818
rect 12835 9766 12849 9818
rect 12873 9766 12887 9818
rect 12887 9766 12899 9818
rect 12899 9766 12929 9818
rect 12953 9766 12963 9818
rect 12963 9766 13009 9818
rect 12713 9764 12769 9766
rect 12793 9764 12849 9766
rect 12873 9764 12929 9766
rect 12953 9764 13009 9766
rect 12438 9560 12494 9616
rect 12053 9274 12109 9276
rect 12133 9274 12189 9276
rect 12213 9274 12269 9276
rect 12293 9274 12349 9276
rect 12053 9222 12099 9274
rect 12099 9222 12109 9274
rect 12133 9222 12163 9274
rect 12163 9222 12175 9274
rect 12175 9222 12189 9274
rect 12213 9222 12227 9274
rect 12227 9222 12239 9274
rect 12239 9222 12269 9274
rect 12293 9222 12303 9274
rect 12303 9222 12349 9274
rect 12053 9220 12109 9222
rect 12133 9220 12189 9222
rect 12213 9220 12269 9222
rect 12293 9220 12349 9222
rect 12622 9152 12678 9208
rect 12990 9424 13046 9480
rect 12713 8730 12769 8732
rect 12793 8730 12849 8732
rect 12873 8730 12929 8732
rect 12953 8730 13009 8732
rect 12713 8678 12759 8730
rect 12759 8678 12769 8730
rect 12793 8678 12823 8730
rect 12823 8678 12835 8730
rect 12835 8678 12849 8730
rect 12873 8678 12887 8730
rect 12887 8678 12899 8730
rect 12899 8678 12929 8730
rect 12953 8678 12963 8730
rect 12963 8678 13009 8730
rect 12713 8676 12769 8678
rect 12793 8676 12849 8678
rect 12873 8676 12929 8678
rect 12953 8676 13009 8678
rect 12530 8608 12586 8664
rect 12053 8186 12109 8188
rect 12133 8186 12189 8188
rect 12213 8186 12269 8188
rect 12293 8186 12349 8188
rect 12053 8134 12099 8186
rect 12099 8134 12109 8186
rect 12133 8134 12163 8186
rect 12163 8134 12175 8186
rect 12175 8134 12189 8186
rect 12213 8134 12227 8186
rect 12227 8134 12239 8186
rect 12239 8134 12269 8186
rect 12293 8134 12303 8186
rect 12303 8134 12349 8186
rect 12053 8132 12109 8134
rect 12133 8132 12189 8134
rect 12213 8132 12269 8134
rect 12293 8132 12349 8134
rect 12530 8084 12586 8120
rect 12530 8064 12532 8084
rect 12532 8064 12584 8084
rect 12584 8064 12586 8084
rect 12254 7928 12310 7984
rect 12530 7928 12586 7984
rect 12254 7792 12310 7848
rect 12162 7520 12218 7576
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 12530 7656 12586 7712
rect 13726 12552 13782 12608
rect 13726 11328 13782 11384
rect 13818 11056 13874 11112
rect 13450 9832 13506 9888
rect 13358 9288 13414 9344
rect 14186 10240 14242 10296
rect 14094 9560 14150 9616
rect 12714 8200 12770 8256
rect 12806 7792 12862 7848
rect 13174 7656 13230 7712
rect 12713 7642 12769 7644
rect 12793 7642 12849 7644
rect 12873 7642 12929 7644
rect 12953 7642 13009 7644
rect 12713 7590 12759 7642
rect 12759 7590 12769 7642
rect 12793 7590 12823 7642
rect 12823 7590 12835 7642
rect 12835 7590 12849 7642
rect 12873 7590 12887 7642
rect 12887 7590 12899 7642
rect 12899 7590 12929 7642
rect 12953 7590 12963 7642
rect 12963 7590 13009 7642
rect 12713 7588 12769 7590
rect 12793 7588 12849 7590
rect 12873 7588 12929 7590
rect 12953 7588 13009 7590
rect 12254 6840 12310 6896
rect 12438 6840 12494 6896
rect 12346 6568 12402 6624
rect 12622 6704 12678 6760
rect 12530 6432 12586 6488
rect 12713 6554 12769 6556
rect 12793 6554 12849 6556
rect 12873 6554 12929 6556
rect 12953 6554 13009 6556
rect 12713 6502 12759 6554
rect 12759 6502 12769 6554
rect 12793 6502 12823 6554
rect 12823 6502 12835 6554
rect 12835 6502 12849 6554
rect 12873 6502 12887 6554
rect 12887 6502 12899 6554
rect 12899 6502 12929 6554
rect 12953 6502 12963 6554
rect 12963 6502 13009 6554
rect 12713 6500 12769 6502
rect 12793 6500 12849 6502
rect 12873 6500 12929 6502
rect 12953 6500 13009 6502
rect 12530 6024 12586 6080
rect 12806 6024 12862 6080
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 12346 3612 12348 3632
rect 12348 3612 12400 3632
rect 12400 3612 12402 3632
rect 12346 3576 12402 3612
rect 11794 3032 11850 3088
rect 12713 5466 12769 5468
rect 12793 5466 12849 5468
rect 12873 5466 12929 5468
rect 12953 5466 13009 5468
rect 12713 5414 12759 5466
rect 12759 5414 12769 5466
rect 12793 5414 12823 5466
rect 12823 5414 12835 5466
rect 12835 5414 12849 5466
rect 12873 5414 12887 5466
rect 12887 5414 12899 5466
rect 12899 5414 12929 5466
rect 12953 5414 12963 5466
rect 12963 5414 13009 5466
rect 12713 5412 12769 5414
rect 12793 5412 12849 5414
rect 12873 5412 12929 5414
rect 12953 5412 13009 5414
rect 12713 4378 12769 4380
rect 12793 4378 12849 4380
rect 12873 4378 12929 4380
rect 12953 4378 13009 4380
rect 12713 4326 12759 4378
rect 12759 4326 12769 4378
rect 12793 4326 12823 4378
rect 12823 4326 12835 4378
rect 12835 4326 12849 4378
rect 12873 4326 12887 4378
rect 12887 4326 12899 4378
rect 12899 4326 12929 4378
rect 12953 4326 12963 4378
rect 12963 4326 13009 4378
rect 12713 4324 12769 4326
rect 12793 4324 12849 4326
rect 12873 4324 12929 4326
rect 12953 4324 13009 4326
rect 12898 4120 12954 4176
rect 12713 3290 12769 3292
rect 12793 3290 12849 3292
rect 12873 3290 12929 3292
rect 12953 3290 13009 3292
rect 12713 3238 12759 3290
rect 12759 3238 12769 3290
rect 12793 3238 12823 3290
rect 12823 3238 12835 3290
rect 12835 3238 12849 3290
rect 12873 3238 12887 3290
rect 12887 3238 12899 3290
rect 12899 3238 12929 3290
rect 12953 3238 12963 3290
rect 12963 3238 13009 3290
rect 12713 3236 12769 3238
rect 12793 3236 12849 3238
rect 12873 3236 12929 3238
rect 12953 3236 13009 3238
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 13450 8880 13506 8936
rect 13818 9016 13874 9072
rect 13818 8336 13874 8392
rect 13726 7268 13782 7304
rect 13726 7248 13728 7268
rect 13728 7248 13780 7268
rect 13780 7248 13782 7268
rect 13450 6976 13506 7032
rect 13358 6840 13414 6896
rect 14002 9424 14058 9480
rect 14554 13096 14610 13152
rect 15566 17856 15622 17912
rect 17958 17720 18014 17776
rect 17152 17434 17208 17436
rect 17232 17434 17288 17436
rect 17312 17434 17368 17436
rect 17392 17434 17448 17436
rect 17152 17382 17198 17434
rect 17198 17382 17208 17434
rect 17232 17382 17262 17434
rect 17262 17382 17274 17434
rect 17274 17382 17288 17434
rect 17312 17382 17326 17434
rect 17326 17382 17338 17434
rect 17338 17382 17368 17434
rect 17392 17382 17402 17434
rect 17402 17382 17448 17434
rect 17152 17380 17208 17382
rect 17232 17380 17288 17382
rect 17312 17380 17368 17382
rect 17392 17380 17448 17382
rect 16492 16890 16548 16892
rect 16572 16890 16628 16892
rect 16652 16890 16708 16892
rect 16732 16890 16788 16892
rect 16492 16838 16538 16890
rect 16538 16838 16548 16890
rect 16572 16838 16602 16890
rect 16602 16838 16614 16890
rect 16614 16838 16628 16890
rect 16652 16838 16666 16890
rect 16666 16838 16678 16890
rect 16678 16838 16708 16890
rect 16732 16838 16742 16890
rect 16742 16838 16788 16890
rect 16492 16836 16548 16838
rect 16572 16836 16628 16838
rect 16652 16836 16708 16838
rect 16732 16836 16788 16838
rect 15750 16652 15806 16688
rect 15750 16632 15752 16652
rect 15752 16632 15804 16652
rect 15804 16632 15806 16652
rect 14922 13640 14978 13696
rect 15566 14456 15622 14512
rect 14462 11636 14464 11656
rect 14464 11636 14516 11656
rect 14516 11636 14518 11656
rect 14462 11600 14518 11636
rect 14370 11056 14426 11112
rect 14922 12144 14978 12200
rect 15106 12552 15162 12608
rect 15290 12416 15346 12472
rect 15014 11192 15070 11248
rect 14922 11092 14924 11112
rect 14924 11092 14976 11112
rect 14976 11092 14978 11112
rect 14922 11056 14978 11092
rect 14462 10376 14518 10432
rect 14370 9424 14426 9480
rect 14370 9324 14372 9344
rect 14372 9324 14424 9344
rect 14424 9324 14426 9344
rect 14370 9288 14426 9324
rect 14002 8744 14058 8800
rect 14002 8336 14058 8392
rect 14002 5888 14058 5944
rect 14186 6160 14242 6216
rect 14738 10512 14794 10568
rect 14646 10412 14648 10432
rect 14648 10412 14700 10432
rect 14700 10412 14702 10432
rect 14646 10376 14702 10412
rect 15198 9016 15254 9072
rect 14738 8336 14794 8392
rect 14646 6840 14702 6896
rect 15014 8200 15070 8256
rect 14554 3576 14610 3632
rect 15106 7656 15162 7712
rect 15566 12708 15622 12744
rect 15566 12688 15568 12708
rect 15568 12688 15620 12708
rect 15620 12688 15622 12708
rect 15566 12552 15622 12608
rect 15474 11736 15530 11792
rect 15658 11736 15714 11792
rect 15658 8880 15714 8936
rect 15566 8064 15622 8120
rect 15474 5616 15530 5672
rect 15934 12300 15990 12336
rect 15934 12280 15936 12300
rect 15936 12280 15988 12300
rect 15988 12280 15990 12300
rect 16492 15802 16548 15804
rect 16572 15802 16628 15804
rect 16652 15802 16708 15804
rect 16732 15802 16788 15804
rect 16492 15750 16538 15802
rect 16538 15750 16548 15802
rect 16572 15750 16602 15802
rect 16602 15750 16614 15802
rect 16614 15750 16628 15802
rect 16652 15750 16666 15802
rect 16666 15750 16678 15802
rect 16678 15750 16708 15802
rect 16732 15750 16742 15802
rect 16742 15750 16788 15802
rect 16492 15748 16548 15750
rect 16572 15748 16628 15750
rect 16652 15748 16708 15750
rect 16732 15748 16788 15750
rect 16492 14714 16548 14716
rect 16572 14714 16628 14716
rect 16652 14714 16708 14716
rect 16732 14714 16788 14716
rect 16492 14662 16538 14714
rect 16538 14662 16548 14714
rect 16572 14662 16602 14714
rect 16602 14662 16614 14714
rect 16614 14662 16628 14714
rect 16652 14662 16666 14714
rect 16666 14662 16678 14714
rect 16678 14662 16708 14714
rect 16732 14662 16742 14714
rect 16742 14662 16788 14714
rect 16492 14660 16548 14662
rect 16572 14660 16628 14662
rect 16652 14660 16708 14662
rect 16732 14660 16788 14662
rect 16492 13626 16548 13628
rect 16572 13626 16628 13628
rect 16652 13626 16708 13628
rect 16732 13626 16788 13628
rect 16492 13574 16538 13626
rect 16538 13574 16548 13626
rect 16572 13574 16602 13626
rect 16602 13574 16614 13626
rect 16614 13574 16628 13626
rect 16652 13574 16666 13626
rect 16666 13574 16678 13626
rect 16678 13574 16708 13626
rect 16732 13574 16742 13626
rect 16742 13574 16788 13626
rect 16492 13572 16548 13574
rect 16572 13572 16628 13574
rect 16652 13572 16708 13574
rect 16732 13572 16788 13574
rect 16026 9424 16082 9480
rect 15382 3984 15438 4040
rect 15474 3732 15530 3768
rect 15474 3712 15476 3732
rect 15476 3712 15528 3732
rect 15528 3712 15530 3732
rect 16486 12688 16542 12744
rect 17774 16496 17830 16552
rect 17152 16346 17208 16348
rect 17232 16346 17288 16348
rect 17312 16346 17368 16348
rect 17392 16346 17448 16348
rect 17152 16294 17198 16346
rect 17198 16294 17208 16346
rect 17232 16294 17262 16346
rect 17262 16294 17274 16346
rect 17274 16294 17288 16346
rect 17312 16294 17326 16346
rect 17326 16294 17338 16346
rect 17338 16294 17368 16346
rect 17392 16294 17402 16346
rect 17402 16294 17448 16346
rect 17152 16292 17208 16294
rect 17232 16292 17288 16294
rect 17312 16292 17368 16294
rect 17392 16292 17448 16294
rect 17152 15258 17208 15260
rect 17232 15258 17288 15260
rect 17312 15258 17368 15260
rect 17392 15258 17448 15260
rect 17152 15206 17198 15258
rect 17198 15206 17208 15258
rect 17232 15206 17262 15258
rect 17262 15206 17274 15258
rect 17274 15206 17288 15258
rect 17312 15206 17326 15258
rect 17326 15206 17338 15258
rect 17338 15206 17368 15258
rect 17392 15206 17402 15258
rect 17402 15206 17448 15258
rect 17152 15204 17208 15206
rect 17232 15204 17288 15206
rect 17312 15204 17368 15206
rect 17392 15204 17448 15206
rect 17498 14320 17554 14376
rect 17152 14170 17208 14172
rect 17232 14170 17288 14172
rect 17312 14170 17368 14172
rect 17392 14170 17448 14172
rect 17152 14118 17198 14170
rect 17198 14118 17208 14170
rect 17232 14118 17262 14170
rect 17262 14118 17274 14170
rect 17274 14118 17288 14170
rect 17312 14118 17326 14170
rect 17326 14118 17338 14170
rect 17338 14118 17368 14170
rect 17392 14118 17402 14170
rect 17402 14118 17448 14170
rect 17152 14116 17208 14118
rect 17232 14116 17288 14118
rect 17312 14116 17368 14118
rect 17392 14116 17448 14118
rect 17152 13082 17208 13084
rect 17232 13082 17288 13084
rect 17312 13082 17368 13084
rect 17392 13082 17448 13084
rect 17152 13030 17198 13082
rect 17198 13030 17208 13082
rect 17232 13030 17262 13082
rect 17262 13030 17274 13082
rect 17274 13030 17288 13082
rect 17312 13030 17326 13082
rect 17326 13030 17338 13082
rect 17338 13030 17368 13082
rect 17392 13030 17402 13082
rect 17402 13030 17448 13082
rect 17152 13028 17208 13030
rect 17232 13028 17288 13030
rect 17312 13028 17368 13030
rect 17392 13028 17448 13030
rect 16492 12538 16548 12540
rect 16572 12538 16628 12540
rect 16652 12538 16708 12540
rect 16732 12538 16788 12540
rect 16492 12486 16538 12538
rect 16538 12486 16548 12538
rect 16572 12486 16602 12538
rect 16602 12486 16614 12538
rect 16614 12486 16628 12538
rect 16652 12486 16666 12538
rect 16666 12486 16678 12538
rect 16678 12486 16708 12538
rect 16732 12486 16742 12538
rect 16742 12486 16788 12538
rect 16492 12484 16548 12486
rect 16572 12484 16628 12486
rect 16652 12484 16708 12486
rect 16732 12484 16788 12486
rect 16394 11736 16450 11792
rect 16492 11450 16548 11452
rect 16572 11450 16628 11452
rect 16652 11450 16708 11452
rect 16732 11450 16788 11452
rect 16492 11398 16538 11450
rect 16538 11398 16548 11450
rect 16572 11398 16602 11450
rect 16602 11398 16614 11450
rect 16614 11398 16628 11450
rect 16652 11398 16666 11450
rect 16666 11398 16678 11450
rect 16678 11398 16708 11450
rect 16732 11398 16742 11450
rect 16742 11398 16788 11450
rect 16492 11396 16548 11398
rect 16572 11396 16628 11398
rect 16652 11396 16708 11398
rect 16732 11396 16788 11398
rect 16578 10648 16634 10704
rect 16946 11192 17002 11248
rect 16854 10920 16910 10976
rect 16762 10804 16818 10840
rect 16762 10784 16764 10804
rect 16764 10784 16816 10804
rect 16816 10784 16818 10804
rect 16394 10512 16450 10568
rect 16492 10362 16548 10364
rect 16572 10362 16628 10364
rect 16652 10362 16708 10364
rect 16732 10362 16788 10364
rect 16492 10310 16538 10362
rect 16538 10310 16548 10362
rect 16572 10310 16602 10362
rect 16602 10310 16614 10362
rect 16614 10310 16628 10362
rect 16652 10310 16666 10362
rect 16666 10310 16678 10362
rect 16678 10310 16708 10362
rect 16732 10310 16742 10362
rect 16742 10310 16788 10362
rect 16492 10308 16548 10310
rect 16572 10308 16628 10310
rect 16652 10308 16708 10310
rect 16732 10308 16788 10310
rect 16486 9560 16542 9616
rect 17222 12844 17278 12880
rect 17222 12824 17224 12844
rect 17224 12824 17276 12844
rect 17276 12824 17278 12844
rect 17152 11994 17208 11996
rect 17232 11994 17288 11996
rect 17312 11994 17368 11996
rect 17392 11994 17448 11996
rect 17152 11942 17198 11994
rect 17198 11942 17208 11994
rect 17232 11942 17262 11994
rect 17262 11942 17274 11994
rect 17274 11942 17288 11994
rect 17312 11942 17326 11994
rect 17326 11942 17338 11994
rect 17338 11942 17368 11994
rect 17392 11942 17402 11994
rect 17402 11942 17448 11994
rect 17152 11940 17208 11942
rect 17232 11940 17288 11942
rect 17312 11940 17368 11942
rect 17392 11940 17448 11942
rect 17152 10906 17208 10908
rect 17232 10906 17288 10908
rect 17312 10906 17368 10908
rect 17392 10906 17448 10908
rect 17152 10854 17198 10906
rect 17198 10854 17208 10906
rect 17232 10854 17262 10906
rect 17262 10854 17274 10906
rect 17274 10854 17288 10906
rect 17312 10854 17326 10906
rect 17326 10854 17338 10906
rect 17338 10854 17368 10906
rect 17392 10854 17402 10906
rect 17402 10854 17448 10906
rect 17152 10852 17208 10854
rect 17232 10852 17288 10854
rect 17312 10852 17368 10854
rect 17392 10852 17448 10854
rect 17038 9968 17094 10024
rect 16946 9696 17002 9752
rect 17152 9818 17208 9820
rect 17232 9818 17288 9820
rect 17312 9818 17368 9820
rect 17392 9818 17448 9820
rect 17152 9766 17198 9818
rect 17198 9766 17208 9818
rect 17232 9766 17262 9818
rect 17262 9766 17274 9818
rect 17274 9766 17288 9818
rect 17312 9766 17326 9818
rect 17326 9766 17338 9818
rect 17338 9766 17368 9818
rect 17392 9766 17402 9818
rect 17402 9766 17448 9818
rect 17152 9764 17208 9766
rect 17232 9764 17288 9766
rect 17312 9764 17368 9766
rect 17392 9764 17448 9766
rect 16492 9274 16548 9276
rect 16572 9274 16628 9276
rect 16652 9274 16708 9276
rect 16732 9274 16788 9276
rect 16492 9222 16538 9274
rect 16538 9222 16548 9274
rect 16572 9222 16602 9274
rect 16602 9222 16614 9274
rect 16614 9222 16628 9274
rect 16652 9222 16666 9274
rect 16666 9222 16678 9274
rect 16678 9222 16708 9274
rect 16732 9222 16742 9274
rect 16742 9222 16788 9274
rect 16492 9220 16548 9222
rect 16572 9220 16628 9222
rect 16652 9220 16708 9222
rect 16732 9220 16788 9222
rect 16946 9424 17002 9480
rect 17314 8880 17370 8936
rect 16854 8336 16910 8392
rect 16492 8186 16548 8188
rect 16572 8186 16628 8188
rect 16652 8186 16708 8188
rect 16732 8186 16788 8188
rect 16492 8134 16538 8186
rect 16538 8134 16548 8186
rect 16572 8134 16602 8186
rect 16602 8134 16614 8186
rect 16614 8134 16628 8186
rect 16652 8134 16666 8186
rect 16666 8134 16678 8186
rect 16678 8134 16708 8186
rect 16732 8134 16742 8186
rect 16742 8134 16788 8186
rect 16492 8132 16548 8134
rect 16572 8132 16628 8134
rect 16652 8132 16708 8134
rect 16732 8132 16788 8134
rect 16394 7656 16450 7712
rect 17152 8730 17208 8732
rect 17232 8730 17288 8732
rect 17312 8730 17368 8732
rect 17392 8730 17448 8732
rect 17152 8678 17198 8730
rect 17198 8678 17208 8730
rect 17232 8678 17262 8730
rect 17262 8678 17274 8730
rect 17274 8678 17288 8730
rect 17312 8678 17326 8730
rect 17326 8678 17338 8730
rect 17338 8678 17368 8730
rect 17392 8678 17402 8730
rect 17402 8678 17448 8730
rect 17152 8676 17208 8678
rect 17232 8676 17288 8678
rect 17312 8676 17368 8678
rect 17392 8676 17448 8678
rect 17038 7928 17094 7984
rect 16394 7520 16450 7576
rect 16210 5616 16266 5672
rect 16210 5208 16266 5264
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 17590 10104 17646 10160
rect 17498 8372 17500 8392
rect 17500 8372 17552 8392
rect 17552 8372 17554 8392
rect 17498 8336 17554 8372
rect 17152 7642 17208 7644
rect 17232 7642 17288 7644
rect 17312 7642 17368 7644
rect 17392 7642 17448 7644
rect 17152 7590 17198 7642
rect 17198 7590 17208 7642
rect 17232 7590 17262 7642
rect 17262 7590 17274 7642
rect 17274 7590 17288 7642
rect 17312 7590 17326 7642
rect 17326 7590 17338 7642
rect 17338 7590 17368 7642
rect 17392 7590 17402 7642
rect 17402 7590 17448 7642
rect 17152 7588 17208 7590
rect 17232 7588 17288 7590
rect 17312 7588 17368 7590
rect 17392 7588 17448 7590
rect 17038 7384 17094 7440
rect 17866 14864 17922 14920
rect 17774 14048 17830 14104
rect 17774 9560 17830 9616
rect 18786 15544 18842 15600
rect 18050 13232 18106 13288
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 17152 6554 17208 6556
rect 17232 6554 17288 6556
rect 17312 6554 17368 6556
rect 17392 6554 17448 6556
rect 17152 6502 17198 6554
rect 17198 6502 17208 6554
rect 17232 6502 17262 6554
rect 17262 6502 17274 6554
rect 17274 6502 17288 6554
rect 17312 6502 17326 6554
rect 17326 6502 17338 6554
rect 17338 6502 17368 6554
rect 17392 6502 17402 6554
rect 17402 6502 17448 6554
rect 17152 6500 17208 6502
rect 17232 6500 17288 6502
rect 17312 6500 17368 6502
rect 17392 6500 17448 6502
rect 16946 6296 17002 6352
rect 17498 6296 17554 6352
rect 16394 5752 16450 5808
rect 17152 5466 17208 5468
rect 17232 5466 17288 5468
rect 17312 5466 17368 5468
rect 17392 5466 17448 5468
rect 17152 5414 17198 5466
rect 17198 5414 17208 5466
rect 17232 5414 17262 5466
rect 17262 5414 17274 5466
rect 17274 5414 17288 5466
rect 17312 5414 17326 5466
rect 17326 5414 17338 5466
rect 17338 5414 17368 5466
rect 17392 5414 17402 5466
rect 17402 5414 17448 5466
rect 17152 5412 17208 5414
rect 17232 5412 17288 5414
rect 17312 5412 17368 5414
rect 17392 5412 17448 5414
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 16854 4684 16910 4720
rect 16854 4664 16856 4684
rect 16856 4664 16908 4684
rect 16908 4664 16910 4684
rect 18050 7792 18106 7848
rect 17774 5072 17830 5128
rect 17152 4378 17208 4380
rect 17232 4378 17288 4380
rect 17312 4378 17368 4380
rect 17392 4378 17448 4380
rect 17152 4326 17198 4378
rect 17198 4326 17208 4378
rect 17232 4326 17262 4378
rect 17262 4326 17274 4378
rect 17274 4326 17288 4378
rect 17312 4326 17326 4378
rect 17326 4326 17338 4378
rect 17338 4326 17368 4378
rect 17392 4326 17402 4378
rect 17402 4326 17448 4378
rect 17152 4324 17208 4326
rect 17232 4324 17288 4326
rect 17312 4324 17368 4326
rect 17392 4324 17448 4326
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 18602 9016 18658 9072
rect 18326 8336 18382 8392
rect 17152 3290 17208 3292
rect 17232 3290 17288 3292
rect 17312 3290 17368 3292
rect 17392 3290 17448 3292
rect 17152 3238 17198 3290
rect 17198 3238 17208 3290
rect 17232 3238 17262 3290
rect 17262 3238 17274 3290
rect 17274 3238 17288 3290
rect 17312 3238 17326 3290
rect 17326 3238 17338 3290
rect 17338 3238 17368 3290
rect 17392 3238 17402 3290
rect 17402 3238 17448 3290
rect 17152 3236 17208 3238
rect 17232 3236 17288 3238
rect 17312 3236 17368 3238
rect 17392 3236 17448 3238
rect 17774 3188 17830 3224
rect 17774 3168 17776 3188
rect 17776 3168 17828 3188
rect 17828 3168 17830 3188
rect 17314 3032 17370 3088
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 19338 8472 19394 8528
rect 12713 2202 12769 2204
rect 12793 2202 12849 2204
rect 12873 2202 12929 2204
rect 12953 2202 13009 2204
rect 12713 2150 12759 2202
rect 12759 2150 12769 2202
rect 12793 2150 12823 2202
rect 12823 2150 12835 2202
rect 12835 2150 12849 2202
rect 12873 2150 12887 2202
rect 12887 2150 12899 2202
rect 12899 2150 12929 2202
rect 12953 2150 12963 2202
rect 12963 2150 13009 2202
rect 12713 2148 12769 2150
rect 12793 2148 12849 2150
rect 12873 2148 12929 2150
rect 12953 2148 13009 2150
rect 17152 2202 17208 2204
rect 17232 2202 17288 2204
rect 17312 2202 17368 2204
rect 17392 2202 17448 2204
rect 17152 2150 17198 2202
rect 17198 2150 17208 2202
rect 17232 2150 17262 2202
rect 17262 2150 17274 2202
rect 17274 2150 17288 2202
rect 17312 2150 17326 2202
rect 17326 2150 17338 2202
rect 17338 2150 17368 2202
rect 17392 2150 17402 2202
rect 17402 2150 17448 2202
rect 17152 2148 17208 2150
rect 17232 2148 17288 2150
rect 17312 2148 17368 2150
rect 17392 2148 17448 2150
<< metal3 >>
rect 0 19818 800 19848
rect 9254 19818 9260 19820
rect 0 19758 9260 19818
rect 0 19728 800 19758
rect 9254 19756 9260 19758
rect 9324 19756 9330 19820
rect 0 19138 800 19168
rect 2865 19138 2931 19141
rect 0 19136 2931 19138
rect 0 19080 2870 19136
rect 2926 19080 2931 19136
rect 0 19078 2931 19080
rect 0 19048 800 19078
rect 2865 19075 2931 19078
rect 0 18458 800 18488
rect 2773 18458 2839 18461
rect 0 18456 2839 18458
rect 0 18400 2778 18456
rect 2834 18400 2839 18456
rect 0 18398 2839 18400
rect 0 18368 800 18398
rect 2773 18395 2839 18398
rect 6729 18186 6795 18189
rect 16982 18186 16988 18188
rect 6729 18184 16988 18186
rect 6729 18128 6734 18184
rect 6790 18128 16988 18184
rect 6729 18126 16988 18128
rect 6729 18123 6795 18126
rect 16982 18124 16988 18126
rect 17052 18124 17058 18188
rect 1342 17988 1348 18052
rect 1412 18050 1418 18052
rect 15377 18050 15443 18053
rect 1412 18048 15443 18050
rect 1412 17992 15382 18048
rect 15438 17992 15443 18048
rect 1412 17990 15443 17992
rect 1412 17988 1418 17990
rect 15377 17987 15443 17990
rect 933 17914 999 17917
rect 15561 17914 15627 17917
rect 933 17912 15627 17914
rect 933 17856 938 17912
rect 994 17856 15566 17912
rect 15622 17856 15627 17912
rect 933 17854 15627 17856
rect 933 17851 999 17854
rect 15561 17851 15627 17854
rect 0 17778 800 17808
rect 2957 17778 3023 17781
rect 0 17776 3023 17778
rect 0 17720 2962 17776
rect 3018 17720 3023 17776
rect 0 17718 3023 17720
rect 0 17688 800 17718
rect 2957 17715 3023 17718
rect 8017 17778 8083 17781
rect 17953 17778 18019 17781
rect 8017 17776 18019 17778
rect 8017 17720 8022 17776
rect 8078 17720 17958 17776
rect 18014 17720 18019 17776
rect 8017 17718 18019 17720
rect 8017 17715 8083 17718
rect 17953 17715 18019 17718
rect 1158 17580 1164 17644
rect 1228 17642 1234 17644
rect 14365 17642 14431 17645
rect 1228 17640 14431 17642
rect 1228 17584 14370 17640
rect 14426 17584 14431 17640
rect 1228 17582 14431 17584
rect 1228 17580 1234 17582
rect 14365 17579 14431 17582
rect 3825 17440 4141 17441
rect 3825 17376 3831 17440
rect 3895 17376 3911 17440
rect 3975 17376 3991 17440
rect 4055 17376 4071 17440
rect 4135 17376 4141 17440
rect 3825 17375 4141 17376
rect 8264 17440 8580 17441
rect 8264 17376 8270 17440
rect 8334 17376 8350 17440
rect 8414 17376 8430 17440
rect 8494 17376 8510 17440
rect 8574 17376 8580 17440
rect 8264 17375 8580 17376
rect 12703 17440 13019 17441
rect 12703 17376 12709 17440
rect 12773 17376 12789 17440
rect 12853 17376 12869 17440
rect 12933 17376 12949 17440
rect 13013 17376 13019 17440
rect 12703 17375 13019 17376
rect 17142 17440 17458 17441
rect 17142 17376 17148 17440
rect 17212 17376 17228 17440
rect 17292 17376 17308 17440
rect 17372 17376 17388 17440
rect 17452 17376 17458 17440
rect 17142 17375 17458 17376
rect 6821 17370 6887 17373
rect 7649 17370 7715 17373
rect 6821 17368 7715 17370
rect 6821 17312 6826 17368
rect 6882 17312 7654 17368
rect 7710 17312 7715 17368
rect 6821 17310 7715 17312
rect 6821 17307 6887 17310
rect 7649 17307 7715 17310
rect 7281 17234 7347 17237
rect 12341 17234 12407 17237
rect 7281 17232 12407 17234
rect 7281 17176 7286 17232
rect 7342 17176 12346 17232
rect 12402 17176 12407 17232
rect 7281 17174 12407 17176
rect 7281 17171 7347 17174
rect 12341 17171 12407 17174
rect 0 17098 800 17128
rect 3049 17098 3115 17101
rect 5073 17098 5139 17101
rect 0 17096 5139 17098
rect 0 17040 3054 17096
rect 3110 17040 5078 17096
rect 5134 17040 5139 17096
rect 0 17038 5139 17040
rect 0 17008 800 17038
rect 3049 17035 3115 17038
rect 5073 17035 5139 17038
rect 12157 17098 12223 17101
rect 17718 17098 17724 17100
rect 12157 17096 17724 17098
rect 12157 17040 12162 17096
rect 12218 17040 17724 17096
rect 12157 17038 17724 17040
rect 12157 17035 12223 17038
rect 17718 17036 17724 17038
rect 17788 17036 17794 17100
rect 9070 16900 9076 16964
rect 9140 16962 9146 16964
rect 9397 16962 9463 16965
rect 9140 16960 9463 16962
rect 9140 16904 9402 16960
rect 9458 16904 9463 16960
rect 9140 16902 9463 16904
rect 9140 16900 9146 16902
rect 9397 16899 9463 16902
rect 3165 16896 3481 16897
rect 3165 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3481 16896
rect 3165 16831 3481 16832
rect 7604 16896 7920 16897
rect 7604 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7920 16896
rect 7604 16831 7920 16832
rect 12043 16896 12359 16897
rect 12043 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12359 16896
rect 12043 16831 12359 16832
rect 16482 16896 16798 16897
rect 16482 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16798 16896
rect 16482 16831 16798 16832
rect 9622 16826 9628 16828
rect 8158 16766 9628 16826
rect 381 16690 447 16693
rect 933 16690 999 16693
rect 381 16688 999 16690
rect 381 16632 386 16688
rect 442 16632 938 16688
rect 994 16632 999 16688
rect 381 16630 999 16632
rect 381 16627 447 16630
rect 933 16627 999 16630
rect 2998 16628 3004 16692
rect 3068 16690 3074 16692
rect 3877 16690 3943 16693
rect 3068 16688 3943 16690
rect 3068 16632 3882 16688
rect 3938 16632 3943 16688
rect 3068 16630 3943 16632
rect 3068 16628 3074 16630
rect 3877 16627 3943 16630
rect 5809 16690 5875 16693
rect 8158 16690 8218 16766
rect 9622 16764 9628 16766
rect 9692 16764 9698 16828
rect 5809 16688 8218 16690
rect 5809 16632 5814 16688
rect 5870 16632 8218 16688
rect 5809 16630 8218 16632
rect 8385 16690 8451 16693
rect 10961 16690 11027 16693
rect 8385 16688 11027 16690
rect 8385 16632 8390 16688
rect 8446 16632 10966 16688
rect 11022 16632 11027 16688
rect 8385 16630 11027 16632
rect 5809 16627 5875 16630
rect 8385 16627 8451 16630
rect 10961 16627 11027 16630
rect 11237 16690 11303 16693
rect 15745 16690 15811 16693
rect 11237 16688 15811 16690
rect 11237 16632 11242 16688
rect 11298 16632 15750 16688
rect 15806 16632 15811 16688
rect 11237 16630 15811 16632
rect 11237 16627 11303 16630
rect 15745 16627 15811 16630
rect 2630 16492 2636 16556
rect 2700 16554 2706 16556
rect 2773 16554 2839 16557
rect 2700 16552 2839 16554
rect 2700 16496 2778 16552
rect 2834 16496 2839 16552
rect 2700 16494 2839 16496
rect 2700 16492 2706 16494
rect 2773 16491 2839 16494
rect 2957 16554 3023 16557
rect 5257 16554 5323 16557
rect 2957 16552 5323 16554
rect 2957 16496 2962 16552
rect 3018 16496 5262 16552
rect 5318 16496 5323 16552
rect 2957 16494 5323 16496
rect 2957 16491 3023 16494
rect 5257 16491 5323 16494
rect 7281 16554 7347 16557
rect 17769 16554 17835 16557
rect 7281 16552 17835 16554
rect 7281 16496 7286 16552
rect 7342 16496 17774 16552
rect 17830 16496 17835 16552
rect 7281 16494 17835 16496
rect 7281 16491 7347 16494
rect 17769 16491 17835 16494
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 3825 16352 4141 16353
rect 3825 16288 3831 16352
rect 3895 16288 3911 16352
rect 3975 16288 3991 16352
rect 4055 16288 4071 16352
rect 4135 16288 4141 16352
rect 3825 16287 4141 16288
rect 8264 16352 8580 16353
rect 8264 16288 8270 16352
rect 8334 16288 8350 16352
rect 8414 16288 8430 16352
rect 8494 16288 8510 16352
rect 8574 16288 8580 16352
rect 8264 16287 8580 16288
rect 12703 16352 13019 16353
rect 12703 16288 12709 16352
rect 12773 16288 12789 16352
rect 12853 16288 12869 16352
rect 12933 16288 12949 16352
rect 13013 16288 13019 16352
rect 12703 16287 13019 16288
rect 17142 16352 17458 16353
rect 17142 16288 17148 16352
rect 17212 16288 17228 16352
rect 17292 16288 17308 16352
rect 17372 16288 17388 16352
rect 17452 16288 17458 16352
rect 17142 16287 17458 16288
rect 4470 16220 4476 16284
rect 4540 16282 4546 16284
rect 7189 16282 7255 16285
rect 4540 16280 7255 16282
rect 4540 16224 7194 16280
rect 7250 16224 7255 16280
rect 4540 16222 7255 16224
rect 4540 16220 4546 16222
rect 7189 16219 7255 16222
rect 9121 16282 9187 16285
rect 9581 16282 9647 16285
rect 9121 16280 9647 16282
rect 9121 16224 9126 16280
rect 9182 16224 9586 16280
rect 9642 16224 9647 16280
rect 9121 16222 9647 16224
rect 9121 16219 9187 16222
rect 9581 16219 9647 16222
rect 9990 16220 9996 16284
rect 10060 16282 10066 16284
rect 12525 16282 12591 16285
rect 10060 16280 12591 16282
rect 10060 16224 12530 16280
rect 12586 16224 12591 16280
rect 10060 16222 12591 16224
rect 10060 16220 10066 16222
rect 12525 16219 12591 16222
rect 2773 16146 2839 16149
rect 3550 16146 3556 16148
rect 2773 16144 3556 16146
rect 2773 16088 2778 16144
rect 2834 16088 3556 16144
rect 2773 16086 3556 16088
rect 2773 16083 2839 16086
rect 3550 16084 3556 16086
rect 3620 16084 3626 16148
rect 4061 16146 4127 16149
rect 12709 16146 12775 16149
rect 4061 16144 12775 16146
rect 4061 16088 4066 16144
rect 4122 16088 12714 16144
rect 12770 16088 12775 16144
rect 4061 16086 12775 16088
rect 4061 16083 4127 16086
rect 12709 16083 12775 16086
rect 2129 16010 2195 16013
rect 8477 16010 8543 16013
rect 2129 16008 8543 16010
rect 2129 15952 2134 16008
rect 2190 15952 8482 16008
rect 8538 15952 8543 16008
rect 2129 15950 8543 15952
rect 2129 15947 2195 15950
rect 8477 15947 8543 15950
rect 9121 16010 9187 16013
rect 14774 16010 14780 16012
rect 9121 16008 14780 16010
rect 9121 15952 9126 16008
rect 9182 15952 14780 16008
rect 9121 15950 14780 15952
rect 9121 15947 9187 15950
rect 14774 15948 14780 15950
rect 14844 15948 14850 16012
rect 841 15874 907 15877
rect 6821 15876 6887 15877
rect 6821 15874 6868 15876
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 6776 15872 6868 15874
rect 6776 15816 6826 15872
rect 6776 15814 6868 15816
rect 6821 15812 6868 15814
rect 6932 15812 6938 15876
rect 8201 15874 8267 15877
rect 8845 15874 8911 15877
rect 8201 15872 8911 15874
rect 8201 15816 8206 15872
rect 8262 15816 8850 15872
rect 8906 15816 8911 15872
rect 8201 15814 8911 15816
rect 6821 15811 6887 15812
rect 8201 15811 8267 15814
rect 8845 15811 8911 15814
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 3165 15808 3481 15809
rect 3165 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3481 15808
rect 3165 15743 3481 15744
rect 7604 15808 7920 15809
rect 7604 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7920 15808
rect 7604 15743 7920 15744
rect 12043 15808 12359 15809
rect 12043 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12359 15808
rect 12043 15743 12359 15744
rect 16482 15808 16798 15809
rect 16482 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16798 15808
rect 16482 15743 16798 15744
rect 0 15648 800 15678
rect 5993 15602 6059 15605
rect 12525 15602 12591 15605
rect 18781 15602 18847 15605
rect 5993 15600 12591 15602
rect 5993 15544 5998 15600
rect 6054 15544 12530 15600
rect 12586 15544 12591 15600
rect 5993 15542 12591 15544
rect 5993 15539 6059 15542
rect 12525 15539 12591 15542
rect 14046 15600 18847 15602
rect 14046 15544 18786 15600
rect 18842 15544 18847 15600
rect 14046 15542 18847 15544
rect 5901 15466 5967 15469
rect 9397 15466 9463 15469
rect 5901 15464 9463 15466
rect 5901 15408 5906 15464
rect 5962 15408 9402 15464
rect 9458 15408 9463 15464
rect 5901 15406 9463 15408
rect 5901 15403 5967 15406
rect 9397 15403 9463 15406
rect 9581 15466 9647 15469
rect 14046 15466 14106 15542
rect 18781 15539 18847 15542
rect 9581 15464 14106 15466
rect 9581 15408 9586 15464
rect 9642 15408 14106 15464
rect 9581 15406 14106 15408
rect 14273 15466 14339 15469
rect 15510 15466 15516 15468
rect 14273 15464 15516 15466
rect 14273 15408 14278 15464
rect 14334 15408 15516 15464
rect 14273 15406 15516 15408
rect 9581 15403 9647 15406
rect 14273 15403 14339 15406
rect 15510 15404 15516 15406
rect 15580 15404 15586 15468
rect 2405 15330 2471 15333
rect 3141 15330 3207 15333
rect 2405 15328 3207 15330
rect 2405 15272 2410 15328
rect 2466 15272 3146 15328
rect 3202 15272 3207 15328
rect 2405 15270 3207 15272
rect 2405 15267 2471 15270
rect 3141 15267 3207 15270
rect 9121 15330 9187 15333
rect 12065 15330 12131 15333
rect 9121 15328 12131 15330
rect 9121 15272 9126 15328
rect 9182 15272 12070 15328
rect 12126 15272 12131 15328
rect 9121 15270 12131 15272
rect 9121 15267 9187 15270
rect 12065 15267 12131 15270
rect 14549 15332 14615 15333
rect 14549 15328 14596 15332
rect 14660 15330 14666 15332
rect 14549 15272 14554 15328
rect 14549 15268 14596 15272
rect 14660 15270 14706 15330
rect 14660 15268 14666 15270
rect 14549 15267 14615 15268
rect 3825 15264 4141 15265
rect 3825 15200 3831 15264
rect 3895 15200 3911 15264
rect 3975 15200 3991 15264
rect 4055 15200 4071 15264
rect 4135 15200 4141 15264
rect 3825 15199 4141 15200
rect 8264 15264 8580 15265
rect 8264 15200 8270 15264
rect 8334 15200 8350 15264
rect 8414 15200 8430 15264
rect 8494 15200 8510 15264
rect 8574 15200 8580 15264
rect 8264 15199 8580 15200
rect 12703 15264 13019 15265
rect 12703 15200 12709 15264
rect 12773 15200 12789 15264
rect 12853 15200 12869 15264
rect 12933 15200 12949 15264
rect 13013 15200 13019 15264
rect 12703 15199 13019 15200
rect 17142 15264 17458 15265
rect 17142 15200 17148 15264
rect 17212 15200 17228 15264
rect 17292 15200 17308 15264
rect 17372 15200 17388 15264
rect 17452 15200 17458 15264
rect 17142 15199 17458 15200
rect 4613 15194 4679 15197
rect 7046 15194 7052 15196
rect 4613 15192 7052 15194
rect 4613 15136 4618 15192
rect 4674 15136 7052 15192
rect 4613 15134 7052 15136
rect 4613 15131 4679 15134
rect 7046 15132 7052 15134
rect 7116 15132 7122 15196
rect 10961 15194 11027 15197
rect 10961 15192 12634 15194
rect 10961 15136 10966 15192
rect 11022 15136 12634 15192
rect 10961 15134 12634 15136
rect 10961 15131 11027 15134
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 2497 15058 2563 15061
rect 5349 15058 5415 15061
rect 2497 15056 5415 15058
rect 2497 15000 2502 15056
rect 2558 15000 5354 15056
rect 5410 15000 5415 15056
rect 2497 14998 5415 15000
rect 2497 14995 2563 14998
rect 5349 14995 5415 14998
rect 5901 15058 5967 15061
rect 12433 15058 12499 15061
rect 5901 15056 12499 15058
rect 5901 15000 5906 15056
rect 5962 15000 12438 15056
rect 12494 15000 12499 15056
rect 5901 14998 12499 15000
rect 12574 15058 12634 15134
rect 17902 15058 17908 15060
rect 12574 14998 17908 15058
rect 5901 14995 5967 14998
rect 12433 14995 12499 14998
rect 17902 14996 17908 14998
rect 17972 14996 17978 15060
rect 4429 14922 4495 14925
rect 7925 14922 7991 14925
rect 4429 14920 7991 14922
rect 4429 14864 4434 14920
rect 4490 14864 7930 14920
rect 7986 14864 7991 14920
rect 4429 14862 7991 14864
rect 4429 14859 4495 14862
rect 7925 14859 7991 14862
rect 9029 14922 9095 14925
rect 14089 14922 14155 14925
rect 17861 14922 17927 14925
rect 9029 14920 14155 14922
rect 9029 14864 9034 14920
rect 9090 14864 14094 14920
rect 14150 14864 14155 14920
rect 9029 14862 14155 14864
rect 9029 14859 9095 14862
rect 14089 14859 14155 14862
rect 16254 14920 17927 14922
rect 16254 14864 17866 14920
rect 17922 14864 17927 14920
rect 16254 14862 17927 14864
rect 8702 14724 8708 14788
rect 8772 14786 8778 14788
rect 12433 14786 12499 14789
rect 16254 14786 16314 14862
rect 17861 14859 17927 14862
rect 8772 14726 11714 14786
rect 8772 14724 8778 14726
rect 3165 14720 3481 14721
rect 3165 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3481 14720
rect 3165 14655 3481 14656
rect 7604 14720 7920 14721
rect 7604 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7920 14720
rect 7604 14655 7920 14656
rect 8201 14650 8267 14653
rect 11462 14650 11468 14652
rect 8201 14648 11468 14650
rect 8201 14592 8206 14648
rect 8262 14592 11468 14648
rect 8201 14590 11468 14592
rect 8201 14587 8267 14590
rect 11462 14588 11468 14590
rect 11532 14588 11538 14652
rect 2221 14514 2287 14517
rect 8109 14514 8175 14517
rect 2221 14512 8175 14514
rect 2221 14456 2226 14512
rect 2282 14456 8114 14512
rect 8170 14456 8175 14512
rect 2221 14454 8175 14456
rect 2221 14451 2287 14454
rect 8109 14451 8175 14454
rect 8477 14514 8543 14517
rect 10041 14514 10107 14517
rect 8477 14512 10107 14514
rect 8477 14456 8482 14512
rect 8538 14456 10046 14512
rect 10102 14456 10107 14512
rect 8477 14454 10107 14456
rect 8477 14451 8543 14454
rect 10041 14451 10107 14454
rect 10225 14514 10291 14517
rect 11094 14514 11100 14516
rect 10225 14512 11100 14514
rect 10225 14456 10230 14512
rect 10286 14456 11100 14512
rect 10225 14454 11100 14456
rect 10225 14451 10291 14454
rect 11094 14452 11100 14454
rect 11164 14452 11170 14516
rect 11654 14514 11714 14726
rect 12433 14784 16314 14786
rect 12433 14728 12438 14784
rect 12494 14728 16314 14784
rect 12433 14726 16314 14728
rect 12433 14723 12499 14726
rect 12043 14720 12359 14721
rect 12043 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12359 14720
rect 12043 14655 12359 14656
rect 16482 14720 16798 14721
rect 16482 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16798 14720
rect 16482 14655 16798 14656
rect 15561 14514 15627 14517
rect 11654 14512 15627 14514
rect 11654 14456 15566 14512
rect 15622 14456 15627 14512
rect 11654 14454 15627 14456
rect 15561 14451 15627 14454
rect 0 14378 800 14408
rect 1209 14378 1275 14381
rect 0 14376 1275 14378
rect 0 14320 1214 14376
rect 1270 14320 1275 14376
rect 0 14318 1275 14320
rect 0 14288 800 14318
rect 1209 14315 1275 14318
rect 1577 14378 1643 14381
rect 17493 14378 17559 14381
rect 1577 14376 17559 14378
rect 1577 14320 1582 14376
rect 1638 14320 17498 14376
rect 17554 14320 17559 14376
rect 1577 14318 17559 14320
rect 1577 14315 1643 14318
rect 17493 14315 17559 14318
rect 4705 14242 4771 14245
rect 8109 14242 8175 14245
rect 10777 14244 10843 14245
rect 4705 14240 8175 14242
rect 4705 14184 4710 14240
rect 4766 14184 8114 14240
rect 8170 14184 8175 14240
rect 4705 14182 8175 14184
rect 4705 14179 4771 14182
rect 8109 14179 8175 14182
rect 10726 14180 10732 14244
rect 10796 14242 10843 14244
rect 10796 14240 10888 14242
rect 10838 14184 10888 14240
rect 10796 14182 10888 14184
rect 10796 14180 10843 14182
rect 10777 14179 10843 14180
rect 3825 14176 4141 14177
rect 3825 14112 3831 14176
rect 3895 14112 3911 14176
rect 3975 14112 3991 14176
rect 4055 14112 4071 14176
rect 4135 14112 4141 14176
rect 3825 14111 4141 14112
rect 8264 14176 8580 14177
rect 8264 14112 8270 14176
rect 8334 14112 8350 14176
rect 8414 14112 8430 14176
rect 8494 14112 8510 14176
rect 8574 14112 8580 14176
rect 8264 14111 8580 14112
rect 12703 14176 13019 14177
rect 12703 14112 12709 14176
rect 12773 14112 12789 14176
rect 12853 14112 12869 14176
rect 12933 14112 12949 14176
rect 13013 14112 13019 14176
rect 12703 14111 13019 14112
rect 17142 14176 17458 14177
rect 17142 14112 17148 14176
rect 17212 14112 17228 14176
rect 17292 14112 17308 14176
rect 17372 14112 17388 14176
rect 17452 14112 17458 14176
rect 17142 14111 17458 14112
rect 790 14044 796 14108
rect 860 14106 866 14108
rect 2681 14106 2747 14109
rect 4337 14108 4403 14109
rect 4286 14106 4292 14108
rect 860 14104 2747 14106
rect 860 14048 2686 14104
rect 2742 14048 2747 14104
rect 860 14046 2747 14048
rect 4246 14046 4292 14106
rect 4356 14104 4403 14108
rect 4398 14048 4403 14104
rect 860 14044 866 14046
rect 2681 14043 2747 14046
rect 4286 14044 4292 14046
rect 4356 14044 4403 14048
rect 4838 14044 4844 14108
rect 4908 14106 4914 14108
rect 7097 14106 7163 14109
rect 4908 14104 7163 14106
rect 4908 14048 7102 14104
rect 7158 14048 7163 14104
rect 4908 14046 7163 14048
rect 4908 14044 4914 14046
rect 4337 14043 4403 14044
rect 7097 14043 7163 14046
rect 17534 14044 17540 14108
rect 17604 14106 17610 14108
rect 17769 14106 17835 14109
rect 17604 14104 17835 14106
rect 17604 14048 17774 14104
rect 17830 14048 17835 14104
rect 17604 14046 17835 14048
rect 17604 14044 17610 14046
rect 17769 14043 17835 14046
rect 1577 13970 1643 13973
rect 8753 13970 8819 13973
rect 1577 13968 8819 13970
rect 1577 13912 1582 13968
rect 1638 13912 8758 13968
rect 8814 13912 8819 13968
rect 1577 13910 8819 13912
rect 1577 13907 1643 13910
rect 8753 13907 8819 13910
rect 9489 13970 9555 13973
rect 10358 13970 10364 13972
rect 9489 13968 10364 13970
rect 9489 13912 9494 13968
rect 9550 13912 10364 13968
rect 9489 13910 10364 13912
rect 9489 13907 9555 13910
rect 10358 13908 10364 13910
rect 10428 13970 10434 13972
rect 12893 13970 12959 13973
rect 10428 13968 12959 13970
rect 10428 13912 12898 13968
rect 12954 13912 12959 13968
rect 10428 13910 12959 13912
rect 10428 13908 10434 13910
rect 12893 13907 12959 13910
rect 974 13772 980 13836
rect 1044 13834 1050 13836
rect 4889 13834 4955 13837
rect 1044 13832 4955 13834
rect 1044 13776 4894 13832
rect 4950 13776 4955 13832
rect 1044 13774 4955 13776
rect 1044 13772 1050 13774
rect 4889 13771 4955 13774
rect 6269 13834 6335 13837
rect 8937 13834 9003 13837
rect 6269 13832 9003 13834
rect 6269 13776 6274 13832
rect 6330 13776 8942 13832
rect 8998 13776 9003 13832
rect 6269 13774 9003 13776
rect 6269 13771 6335 13774
rect 8937 13771 9003 13774
rect 11654 13774 12588 13834
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 5441 13698 5507 13701
rect 6913 13698 6979 13701
rect 5441 13696 6979 13698
rect 5441 13640 5446 13696
rect 5502 13640 6918 13696
rect 6974 13640 6979 13696
rect 5441 13638 6979 13640
rect 5441 13635 5507 13638
rect 6913 13635 6979 13638
rect 8017 13698 8083 13701
rect 11654 13698 11714 13774
rect 8017 13696 11714 13698
rect 8017 13640 8022 13696
rect 8078 13640 11714 13696
rect 8017 13638 11714 13640
rect 11789 13700 11855 13701
rect 11789 13696 11836 13700
rect 11900 13698 11906 13700
rect 12528 13698 12588 13774
rect 13302 13772 13308 13836
rect 13372 13834 13378 13836
rect 13721 13834 13787 13837
rect 13372 13832 13787 13834
rect 13372 13776 13726 13832
rect 13782 13776 13787 13832
rect 13372 13774 13787 13776
rect 13372 13772 13378 13774
rect 13721 13771 13787 13774
rect 14038 13698 14044 13700
rect 11789 13640 11794 13696
rect 8017 13635 8083 13638
rect 11789 13636 11836 13640
rect 11900 13638 11946 13698
rect 12528 13638 14044 13698
rect 11900 13636 11906 13638
rect 14038 13636 14044 13638
rect 14108 13698 14114 13700
rect 14181 13698 14247 13701
rect 14108 13696 14247 13698
rect 14108 13640 14186 13696
rect 14242 13640 14247 13696
rect 14108 13638 14247 13640
rect 14108 13636 14114 13638
rect 11789 13635 11855 13636
rect 14181 13635 14247 13638
rect 14917 13698 14983 13701
rect 15142 13698 15148 13700
rect 14917 13696 15148 13698
rect 14917 13640 14922 13696
rect 14978 13640 15148 13696
rect 14917 13638 15148 13640
rect 14917 13635 14983 13638
rect 15142 13636 15148 13638
rect 15212 13636 15218 13700
rect 3165 13632 3481 13633
rect 3165 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3481 13632
rect 3165 13567 3481 13568
rect 7604 13632 7920 13633
rect 7604 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7920 13632
rect 7604 13567 7920 13568
rect 12043 13632 12359 13633
rect 12043 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12359 13632
rect 12043 13567 12359 13568
rect 16482 13632 16798 13633
rect 16482 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16798 13632
rect 16482 13567 16798 13568
rect 3969 13562 4035 13565
rect 5257 13562 5323 13565
rect 5441 13562 5507 13565
rect 3969 13560 5507 13562
rect 3969 13504 3974 13560
rect 4030 13504 5262 13560
rect 5318 13504 5446 13560
rect 5502 13504 5507 13560
rect 3969 13502 5507 13504
rect 3969 13499 4035 13502
rect 5257 13499 5323 13502
rect 5441 13499 5507 13502
rect 6177 13562 6243 13565
rect 6494 13562 6500 13564
rect 6177 13560 6500 13562
rect 6177 13504 6182 13560
rect 6238 13504 6500 13560
rect 6177 13502 6500 13504
rect 6177 13499 6243 13502
rect 6494 13500 6500 13502
rect 6564 13500 6570 13564
rect 13813 13426 13879 13429
rect 2730 13424 13879 13426
rect 2730 13368 13818 13424
rect 13874 13368 13879 13424
rect 2730 13366 13879 13368
rect 0 13018 800 13048
rect 1945 13018 2011 13021
rect 0 13016 2011 13018
rect 0 12960 1950 13016
rect 2006 12960 2011 13016
rect 0 12958 2011 12960
rect 0 12928 800 12958
rect 1945 12955 2011 12958
rect 1209 12882 1275 12885
rect 2730 12882 2790 13366
rect 13813 13363 13879 13366
rect 3601 13290 3667 13293
rect 9438 13290 9444 13292
rect 3601 13288 9444 13290
rect 3601 13232 3606 13288
rect 3662 13232 9444 13288
rect 3601 13230 9444 13232
rect 3601 13227 3667 13230
rect 9438 13228 9444 13230
rect 9508 13228 9514 13292
rect 11237 13290 11303 13293
rect 12065 13290 12131 13293
rect 18045 13290 18111 13293
rect 9630 13288 18111 13290
rect 9630 13232 11242 13288
rect 11298 13232 12070 13288
rect 12126 13232 18050 13288
rect 18106 13232 18111 13288
rect 9630 13230 18111 13232
rect 5073 13154 5139 13157
rect 7230 13154 7236 13156
rect 5073 13152 7236 13154
rect 5073 13096 5078 13152
rect 5134 13096 7236 13152
rect 5073 13094 7236 13096
rect 5073 13091 5139 13094
rect 7230 13092 7236 13094
rect 7300 13092 7306 13156
rect 9213 13154 9279 13157
rect 9630 13154 9690 13230
rect 11237 13227 11303 13230
rect 12065 13227 12131 13230
rect 18045 13227 18111 13230
rect 9213 13152 9690 13154
rect 9213 13096 9218 13152
rect 9274 13096 9690 13152
rect 9213 13094 9690 13096
rect 9213 13091 9279 13094
rect 9806 13092 9812 13156
rect 9876 13154 9882 13156
rect 10133 13154 10199 13157
rect 9876 13152 10199 13154
rect 9876 13096 10138 13152
rect 10194 13096 10199 13152
rect 9876 13094 10199 13096
rect 9876 13092 9882 13094
rect 10133 13091 10199 13094
rect 13905 13154 13971 13157
rect 14089 13154 14155 13157
rect 14549 13154 14615 13157
rect 13905 13152 14615 13154
rect 13905 13096 13910 13152
rect 13966 13096 14094 13152
rect 14150 13096 14554 13152
rect 14610 13096 14615 13152
rect 13905 13094 14615 13096
rect 13905 13091 13971 13094
rect 14089 13091 14155 13094
rect 14549 13091 14615 13094
rect 3825 13088 4141 13089
rect 3825 13024 3831 13088
rect 3895 13024 3911 13088
rect 3975 13024 3991 13088
rect 4055 13024 4071 13088
rect 4135 13024 4141 13088
rect 3825 13023 4141 13024
rect 8264 13088 8580 13089
rect 8264 13024 8270 13088
rect 8334 13024 8350 13088
rect 8414 13024 8430 13088
rect 8494 13024 8510 13088
rect 8574 13024 8580 13088
rect 8264 13023 8580 13024
rect 12703 13088 13019 13089
rect 12703 13024 12709 13088
rect 12773 13024 12789 13088
rect 12853 13024 12869 13088
rect 12933 13024 12949 13088
rect 13013 13024 13019 13088
rect 12703 13023 13019 13024
rect 17142 13088 17458 13089
rect 17142 13024 17148 13088
rect 17212 13024 17228 13088
rect 17292 13024 17308 13088
rect 17372 13024 17388 13088
rect 17452 13024 17458 13088
rect 17142 13023 17458 13024
rect 4245 13018 4311 13021
rect 7557 13018 7623 13021
rect 4245 13016 7623 13018
rect 4245 12960 4250 13016
rect 4306 12960 7562 13016
rect 7618 12960 7623 13016
rect 4245 12958 7623 12960
rect 4245 12955 4311 12958
rect 7557 12955 7623 12958
rect 8753 13018 8819 13021
rect 8753 13016 12634 13018
rect 8753 12960 8758 13016
rect 8814 12960 12634 13016
rect 8753 12958 12634 12960
rect 8753 12955 8819 12958
rect 11789 12882 11855 12885
rect 1209 12880 2790 12882
rect 1209 12824 1214 12880
rect 1270 12824 2790 12880
rect 1209 12822 2790 12824
rect 5950 12880 11855 12882
rect 5950 12824 11794 12880
rect 11850 12824 11855 12880
rect 5950 12822 11855 12824
rect 12574 12882 12634 12958
rect 17217 12882 17283 12885
rect 12574 12880 17283 12882
rect 12574 12824 17222 12880
rect 17278 12824 17283 12880
rect 12574 12822 17283 12824
rect 1209 12819 1275 12822
rect 3550 12684 3556 12748
rect 3620 12746 3626 12748
rect 5950 12746 6010 12822
rect 11789 12819 11855 12822
rect 17217 12819 17283 12822
rect 8477 12746 8543 12749
rect 12249 12746 12315 12749
rect 3620 12686 6010 12746
rect 6318 12686 8080 12746
rect 3620 12684 3626 12686
rect 5165 12610 5231 12613
rect 3558 12608 5231 12610
rect 3558 12552 5170 12608
rect 5226 12552 5231 12608
rect 3558 12550 5231 12552
rect 3165 12544 3481 12545
rect 3165 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3481 12544
rect 3165 12479 3481 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 1577 12338 1643 12341
rect 3558 12338 3618 12550
rect 5165 12547 5231 12550
rect 6085 12612 6151 12613
rect 6085 12608 6132 12612
rect 6196 12610 6202 12612
rect 6085 12552 6090 12608
rect 6085 12548 6132 12552
rect 6196 12550 6242 12610
rect 6196 12548 6202 12550
rect 6085 12547 6151 12548
rect 3693 12474 3759 12477
rect 5022 12474 5028 12476
rect 3693 12472 5028 12474
rect 3693 12416 3698 12472
rect 3754 12416 5028 12472
rect 3693 12414 5028 12416
rect 3693 12411 3759 12414
rect 5022 12412 5028 12414
rect 5092 12474 5098 12476
rect 6318 12474 6378 12686
rect 8020 12610 8080 12686
rect 8477 12744 12315 12746
rect 8477 12688 8482 12744
rect 8538 12688 12254 12744
rect 12310 12688 12315 12744
rect 8477 12686 12315 12688
rect 8477 12683 8543 12686
rect 12249 12683 12315 12686
rect 12801 12746 12867 12749
rect 15561 12746 15627 12749
rect 16481 12746 16547 12749
rect 12801 12744 15627 12746
rect 12801 12688 12806 12744
rect 12862 12688 15566 12744
rect 15622 12688 15627 12744
rect 12801 12686 15627 12688
rect 12801 12683 12867 12686
rect 15561 12683 15627 12686
rect 15702 12744 16547 12746
rect 15702 12688 16486 12744
rect 16542 12688 16547 12744
rect 15702 12686 16547 12688
rect 9213 12610 9279 12613
rect 9806 12610 9812 12612
rect 8020 12608 9279 12610
rect 8020 12552 9218 12608
rect 9274 12552 9279 12608
rect 8020 12550 9279 12552
rect 9213 12547 9279 12550
rect 9630 12550 9812 12610
rect 7604 12544 7920 12545
rect 7604 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7920 12544
rect 7604 12479 7920 12480
rect 5092 12414 6378 12474
rect 9630 12477 9690 12550
rect 9806 12548 9812 12550
rect 9876 12548 9882 12612
rect 10409 12610 10475 12613
rect 11329 12610 11395 12613
rect 10409 12608 11395 12610
rect 10409 12552 10414 12608
rect 10470 12552 11334 12608
rect 11390 12552 11395 12608
rect 10409 12550 11395 12552
rect 10409 12547 10475 12550
rect 11329 12547 11395 12550
rect 13721 12610 13787 12613
rect 15101 12610 15167 12613
rect 13721 12608 15167 12610
rect 13721 12552 13726 12608
rect 13782 12552 15106 12608
rect 15162 12552 15167 12608
rect 13721 12550 15167 12552
rect 13721 12547 13787 12550
rect 15101 12547 15167 12550
rect 15561 12610 15627 12613
rect 15702 12610 15762 12686
rect 16481 12683 16547 12686
rect 15561 12608 15762 12610
rect 15561 12552 15566 12608
rect 15622 12552 15762 12608
rect 15561 12550 15762 12552
rect 15561 12547 15627 12550
rect 12043 12544 12359 12545
rect 12043 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12359 12544
rect 12043 12479 12359 12480
rect 16482 12544 16798 12545
rect 16482 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16798 12544
rect 16482 12479 16798 12480
rect 9630 12472 9739 12477
rect 9630 12416 9678 12472
rect 9734 12416 9739 12472
rect 9630 12414 9739 12416
rect 5092 12412 5098 12414
rect 9673 12411 9739 12414
rect 13077 12474 13143 12477
rect 15285 12474 15351 12477
rect 13077 12472 15351 12474
rect 13077 12416 13082 12472
rect 13138 12416 15290 12472
rect 15346 12416 15351 12472
rect 13077 12414 15351 12416
rect 13077 12411 13143 12414
rect 15285 12411 15351 12414
rect 4245 12340 4311 12341
rect 4245 12338 4292 12340
rect 1577 12336 3618 12338
rect 1577 12280 1582 12336
rect 1638 12280 3618 12336
rect 1577 12278 3618 12280
rect 4200 12336 4292 12338
rect 4200 12280 4250 12336
rect 4200 12278 4292 12280
rect 1577 12275 1643 12278
rect 4245 12276 4292 12278
rect 4356 12276 4362 12340
rect 8109 12338 8175 12341
rect 8702 12338 8708 12340
rect 8109 12336 8708 12338
rect 8109 12280 8114 12336
rect 8170 12280 8708 12336
rect 8109 12278 8708 12280
rect 4245 12275 4311 12276
rect 8109 12275 8175 12278
rect 8702 12276 8708 12278
rect 8772 12276 8778 12340
rect 9806 12276 9812 12340
rect 9876 12338 9882 12340
rect 10409 12338 10475 12341
rect 9876 12336 10475 12338
rect 9876 12280 10414 12336
rect 10470 12280 10475 12336
rect 9876 12278 10475 12280
rect 9876 12276 9882 12278
rect 10409 12275 10475 12278
rect 12433 12338 12499 12341
rect 15929 12338 15995 12341
rect 12433 12336 15995 12338
rect 12433 12280 12438 12336
rect 12494 12280 15934 12336
rect 15990 12280 15995 12336
rect 12433 12278 15995 12280
rect 12433 12275 12499 12278
rect 15929 12275 15995 12278
rect 1209 12202 1275 12205
rect 4889 12202 4955 12205
rect 11053 12202 11119 12205
rect 1209 12200 11119 12202
rect 1209 12144 1214 12200
rect 1270 12144 4894 12200
rect 4950 12144 11058 12200
rect 11114 12144 11119 12200
rect 1209 12142 11119 12144
rect 1209 12139 1275 12142
rect 4889 12139 4955 12142
rect 11053 12139 11119 12142
rect 11646 12140 11652 12204
rect 11716 12202 11722 12204
rect 14917 12202 14983 12205
rect 11716 12200 14983 12202
rect 11716 12144 14922 12200
rect 14978 12144 14983 12200
rect 11716 12142 14983 12144
rect 11716 12140 11722 12142
rect 14917 12139 14983 12142
rect 5441 12066 5507 12069
rect 6678 12066 6684 12068
rect 5441 12064 6684 12066
rect 5441 12008 5446 12064
rect 5502 12008 6684 12064
rect 5441 12006 6684 12008
rect 5441 12003 5507 12006
rect 6678 12004 6684 12006
rect 6748 12004 6754 12068
rect 6821 12066 6887 12069
rect 8017 12066 8083 12069
rect 6821 12064 8083 12066
rect 6821 12008 6826 12064
rect 6882 12008 8022 12064
rect 8078 12008 8083 12064
rect 6821 12006 8083 12008
rect 6821 12003 6887 12006
rect 8017 12003 8083 12006
rect 3825 12000 4141 12001
rect 3825 11936 3831 12000
rect 3895 11936 3911 12000
rect 3975 11936 3991 12000
rect 4055 11936 4071 12000
rect 4135 11936 4141 12000
rect 3825 11935 4141 11936
rect 8264 12000 8580 12001
rect 8264 11936 8270 12000
rect 8334 11936 8350 12000
rect 8414 11936 8430 12000
rect 8494 11936 8510 12000
rect 8574 11936 8580 12000
rect 8264 11935 8580 11936
rect 12703 12000 13019 12001
rect 12703 11936 12709 12000
rect 12773 11936 12789 12000
rect 12853 11936 12869 12000
rect 12933 11936 12949 12000
rect 13013 11936 13019 12000
rect 12703 11935 13019 11936
rect 17142 12000 17458 12001
rect 17142 11936 17148 12000
rect 17212 11936 17228 12000
rect 17292 11936 17308 12000
rect 17372 11936 17388 12000
rect 17452 11936 17458 12000
rect 17142 11935 17458 11936
rect 7414 11868 7420 11932
rect 7484 11930 7490 11932
rect 7741 11930 7807 11933
rect 7484 11928 7807 11930
rect 7484 11872 7746 11928
rect 7802 11872 7807 11928
rect 7484 11870 7807 11872
rect 7484 11868 7490 11870
rect 7741 11867 7807 11870
rect 9213 11930 9279 11933
rect 9806 11930 9812 11932
rect 9213 11928 9812 11930
rect 9213 11872 9218 11928
rect 9274 11872 9812 11928
rect 9213 11870 9812 11872
rect 9213 11867 9279 11870
rect 9806 11868 9812 11870
rect 9876 11868 9882 11932
rect 10174 11868 10180 11932
rect 10244 11930 10250 11932
rect 12433 11930 12499 11933
rect 10244 11928 12499 11930
rect 10244 11872 12438 11928
rect 12494 11872 12499 11928
rect 10244 11870 12499 11872
rect 10244 11868 10250 11870
rect 12433 11867 12499 11870
rect 13445 11930 13511 11933
rect 13670 11930 13676 11932
rect 13445 11928 13676 11930
rect 13445 11872 13450 11928
rect 13506 11872 13676 11928
rect 13445 11870 13676 11872
rect 13445 11867 13511 11870
rect 13670 11868 13676 11870
rect 13740 11868 13746 11932
rect 4429 11794 4495 11797
rect 11329 11794 11395 11797
rect 4429 11792 11395 11794
rect 4429 11736 4434 11792
rect 4490 11736 11334 11792
rect 11390 11736 11395 11792
rect 4429 11734 11395 11736
rect 4429 11731 4495 11734
rect 11329 11731 11395 11734
rect 12893 11794 12959 11797
rect 15469 11794 15535 11797
rect 12893 11792 15535 11794
rect 12893 11736 12898 11792
rect 12954 11736 15474 11792
rect 15530 11736 15535 11792
rect 12893 11734 15535 11736
rect 12893 11731 12959 11734
rect 15469 11731 15535 11734
rect 15653 11794 15719 11797
rect 16389 11794 16455 11797
rect 15653 11792 16455 11794
rect 15653 11736 15658 11792
rect 15714 11736 16394 11792
rect 16450 11736 16455 11792
rect 15653 11734 16455 11736
rect 15653 11731 15719 11734
rect 16389 11731 16455 11734
rect 0 11658 800 11688
rect 1577 11658 1643 11661
rect 0 11656 1643 11658
rect 0 11600 1582 11656
rect 1638 11600 1643 11656
rect 0 11598 1643 11600
rect 0 11568 800 11598
rect 1577 11595 1643 11598
rect 4613 11658 4679 11661
rect 4613 11656 8218 11658
rect 4613 11600 4618 11656
rect 4674 11600 8218 11656
rect 4613 11598 8218 11600
rect 4613 11595 4679 11598
rect 8158 11522 8218 11598
rect 8886 11596 8892 11660
rect 8956 11658 8962 11660
rect 9581 11658 9647 11661
rect 8956 11656 9647 11658
rect 8956 11600 9586 11656
rect 9642 11600 9647 11656
rect 8956 11598 9647 11600
rect 8956 11596 8962 11598
rect 9581 11595 9647 11598
rect 10041 11658 10107 11661
rect 14457 11658 14523 11661
rect 10041 11656 14523 11658
rect 10041 11600 10046 11656
rect 10102 11600 14462 11656
rect 14518 11600 14523 11656
rect 10041 11598 14523 11600
rect 10041 11595 10107 11598
rect 14457 11595 14523 11598
rect 10317 11522 10383 11525
rect 10726 11522 10732 11524
rect 8158 11520 10732 11522
rect 8158 11464 10322 11520
rect 10378 11464 10732 11520
rect 8158 11462 10732 11464
rect 10317 11459 10383 11462
rect 10726 11460 10732 11462
rect 10796 11460 10802 11524
rect 12433 11522 12499 11525
rect 13353 11522 13419 11525
rect 12433 11520 13419 11522
rect 12433 11464 12438 11520
rect 12494 11464 13358 11520
rect 13414 11464 13419 11520
rect 12433 11462 13419 11464
rect 12433 11459 12499 11462
rect 13353 11459 13419 11462
rect 3165 11456 3481 11457
rect 3165 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3481 11456
rect 3165 11391 3481 11392
rect 7604 11456 7920 11457
rect 7604 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7920 11456
rect 7604 11391 7920 11392
rect 12043 11456 12359 11457
rect 12043 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12359 11456
rect 12043 11391 12359 11392
rect 16482 11456 16798 11457
rect 16482 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16798 11456
rect 16482 11391 16798 11392
rect 5165 11386 5231 11389
rect 8385 11386 8451 11389
rect 10501 11388 10567 11389
rect 10501 11386 10548 11388
rect 5165 11384 5274 11386
rect 5165 11328 5170 11384
rect 5226 11328 5274 11384
rect 5165 11323 5274 11328
rect 8385 11384 10548 11386
rect 8385 11328 8390 11384
rect 8446 11328 10506 11384
rect 8385 11326 10548 11328
rect 8385 11323 8451 11326
rect 10501 11324 10548 11326
rect 10612 11324 10618 11388
rect 13721 11386 13787 11389
rect 13721 11384 16314 11386
rect 13721 11328 13726 11384
rect 13782 11328 16314 11384
rect 13721 11326 16314 11328
rect 10501 11323 10567 11324
rect 13721 11323 13787 11326
rect 2313 11250 2379 11253
rect 4838 11250 4844 11252
rect 2313 11248 4844 11250
rect 2313 11192 2318 11248
rect 2374 11192 4844 11248
rect 2313 11190 4844 11192
rect 2313 11187 2379 11190
rect 4838 11188 4844 11190
rect 4908 11188 4914 11252
rect 5214 11250 5274 11323
rect 15009 11250 15075 11253
rect 5214 11248 15075 11250
rect 5214 11192 15014 11248
rect 15070 11192 15075 11248
rect 5214 11190 15075 11192
rect 16254 11250 16314 11326
rect 16941 11250 17007 11253
rect 16254 11248 17007 11250
rect 16254 11192 16946 11248
rect 17002 11192 17007 11248
rect 16254 11190 17007 11192
rect 15009 11187 15075 11190
rect 16941 11187 17007 11190
rect 4705 11114 4771 11117
rect 7281 11114 7347 11117
rect 13353 11114 13419 11117
rect 13813 11114 13879 11117
rect 14365 11116 14431 11117
rect 14917 11116 14983 11117
rect 14365 11114 14412 11116
rect 4705 11112 7114 11114
rect 4705 11056 4710 11112
rect 4766 11056 7114 11112
rect 4705 11054 7114 11056
rect 4705 11051 4771 11054
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 5809 10978 5875 10981
rect 6729 10978 6795 10981
rect 5809 10976 6795 10978
rect 5809 10920 5814 10976
rect 5870 10920 6734 10976
rect 6790 10920 6795 10976
rect 5809 10918 6795 10920
rect 7054 10978 7114 11054
rect 7281 11112 13186 11114
rect 7281 11056 7286 11112
rect 7342 11056 13186 11112
rect 7281 11054 13186 11056
rect 7281 11051 7347 11054
rect 7649 10978 7715 10981
rect 7054 10976 7715 10978
rect 7054 10920 7654 10976
rect 7710 10920 7715 10976
rect 7054 10918 7715 10920
rect 5809 10915 5875 10918
rect 6729 10915 6795 10918
rect 7649 10915 7715 10918
rect 8702 10916 8708 10980
rect 8772 10978 8778 10980
rect 13126 10978 13186 11054
rect 13353 11112 13879 11114
rect 13353 11056 13358 11112
rect 13414 11056 13818 11112
rect 13874 11056 13879 11112
rect 13353 11054 13879 11056
rect 14320 11112 14412 11114
rect 14320 11056 14370 11112
rect 14320 11054 14412 11056
rect 13353 11051 13419 11054
rect 13813 11051 13879 11054
rect 14365 11052 14412 11054
rect 14476 11052 14482 11116
rect 14917 11112 14964 11116
rect 15028 11114 15034 11116
rect 14917 11056 14922 11112
rect 14917 11052 14964 11056
rect 15028 11054 15074 11114
rect 15028 11052 15034 11054
rect 14365 11051 14431 11052
rect 14917 11051 14983 11052
rect 16849 10978 16915 10981
rect 8772 10918 12634 10978
rect 13126 10976 16915 10978
rect 13126 10920 16854 10976
rect 16910 10920 16915 10976
rect 13126 10918 16915 10920
rect 8772 10916 8778 10918
rect 3825 10912 4141 10913
rect 3825 10848 3831 10912
rect 3895 10848 3911 10912
rect 3975 10848 3991 10912
rect 4055 10848 4071 10912
rect 4135 10848 4141 10912
rect 3825 10847 4141 10848
rect 8264 10912 8580 10913
rect 8264 10848 8270 10912
rect 8334 10848 8350 10912
rect 8414 10848 8430 10912
rect 8494 10848 8510 10912
rect 8574 10848 8580 10912
rect 8264 10847 8580 10848
rect 4521 10842 4587 10845
rect 5165 10842 5231 10845
rect 4521 10840 5231 10842
rect 4521 10784 4526 10840
rect 4582 10784 5170 10840
rect 5226 10784 5231 10840
rect 4521 10782 5231 10784
rect 4521 10779 4587 10782
rect 5165 10779 5231 10782
rect 5533 10842 5599 10845
rect 7741 10842 7807 10845
rect 12433 10842 12499 10845
rect 5533 10840 7807 10842
rect 5533 10784 5538 10840
rect 5594 10784 7746 10840
rect 7802 10784 7807 10840
rect 5533 10782 7807 10784
rect 5533 10779 5599 10782
rect 7741 10779 7807 10782
rect 8710 10840 12499 10842
rect 8710 10784 12438 10840
rect 12494 10784 12499 10840
rect 8710 10782 12499 10784
rect 3325 10706 3391 10709
rect 5390 10706 5396 10708
rect 3325 10704 5396 10706
rect 3325 10648 3330 10704
rect 3386 10648 5396 10704
rect 3325 10646 5396 10648
rect 3325 10643 3391 10646
rect 5390 10644 5396 10646
rect 5460 10644 5466 10708
rect 6637 10706 6703 10709
rect 8569 10706 8635 10709
rect 6637 10704 8635 10706
rect 6637 10648 6642 10704
rect 6698 10648 8574 10704
rect 8630 10648 8635 10704
rect 6637 10646 8635 10648
rect 6637 10643 6703 10646
rect 8569 10643 8635 10646
rect 1577 10570 1643 10573
rect 4286 10570 4292 10572
rect 1577 10568 4292 10570
rect 1577 10512 1582 10568
rect 1638 10512 4292 10568
rect 1577 10510 4292 10512
rect 1577 10507 1643 10510
rect 4286 10508 4292 10510
rect 4356 10570 4362 10572
rect 8710 10570 8770 10782
rect 12433 10779 12499 10782
rect 9029 10708 9095 10709
rect 9029 10706 9076 10708
rect 8984 10704 9076 10706
rect 8984 10648 9034 10704
rect 8984 10646 9076 10648
rect 9029 10644 9076 10646
rect 9140 10644 9146 10708
rect 9397 10706 9463 10709
rect 10225 10706 10291 10709
rect 10358 10706 10364 10708
rect 9397 10704 10364 10706
rect 9397 10648 9402 10704
rect 9458 10648 10230 10704
rect 10286 10648 10364 10704
rect 9397 10646 10364 10648
rect 9029 10643 9095 10644
rect 9397 10643 9463 10646
rect 10225 10643 10291 10646
rect 10358 10644 10364 10646
rect 10428 10644 10434 10708
rect 11094 10644 11100 10708
rect 11164 10706 11170 10708
rect 11237 10706 11303 10709
rect 11164 10704 11303 10706
rect 11164 10648 11242 10704
rect 11298 10648 11303 10704
rect 11164 10646 11303 10648
rect 11164 10644 11170 10646
rect 11237 10643 11303 10646
rect 11830 10644 11836 10708
rect 11900 10706 11906 10708
rect 12433 10706 12499 10709
rect 11900 10704 12499 10706
rect 11900 10648 12438 10704
rect 12494 10648 12499 10704
rect 11900 10646 12499 10648
rect 12574 10706 12634 10918
rect 16849 10915 16915 10918
rect 12703 10912 13019 10913
rect 12703 10848 12709 10912
rect 12773 10848 12789 10912
rect 12853 10848 12869 10912
rect 12933 10848 12949 10912
rect 13013 10848 13019 10912
rect 12703 10847 13019 10848
rect 17142 10912 17458 10913
rect 17142 10848 17148 10912
rect 17212 10848 17228 10912
rect 17292 10848 17308 10912
rect 17372 10848 17388 10912
rect 17452 10848 17458 10912
rect 17142 10847 17458 10848
rect 13261 10842 13327 10845
rect 16757 10842 16823 10845
rect 13261 10840 16823 10842
rect 13261 10784 13266 10840
rect 13322 10784 16762 10840
rect 16818 10784 16823 10840
rect 13261 10782 16823 10784
rect 13261 10779 13327 10782
rect 16757 10779 16823 10782
rect 16573 10706 16639 10709
rect 12574 10704 16639 10706
rect 12574 10648 16578 10704
rect 16634 10648 16639 10704
rect 12574 10646 16639 10648
rect 11900 10644 11906 10646
rect 12433 10643 12499 10646
rect 16573 10643 16639 10646
rect 10041 10570 10107 10573
rect 4356 10510 8770 10570
rect 8848 10568 10107 10570
rect 8848 10512 10046 10568
rect 10102 10512 10107 10568
rect 8848 10510 10107 10512
rect 4356 10508 4362 10510
rect 4061 10434 4127 10437
rect 4470 10434 4476 10436
rect 4061 10432 4476 10434
rect 4061 10376 4066 10432
rect 4122 10376 4476 10432
rect 4061 10374 4476 10376
rect 4061 10371 4127 10374
rect 4470 10372 4476 10374
rect 4540 10372 4546 10436
rect 6453 10434 6519 10437
rect 6862 10434 6868 10436
rect 6453 10432 6868 10434
rect 6453 10376 6458 10432
rect 6514 10376 6868 10432
rect 6453 10374 6868 10376
rect 6453 10371 6519 10374
rect 6862 10372 6868 10374
rect 6932 10372 6938 10436
rect 8477 10434 8543 10437
rect 8702 10434 8708 10436
rect 8477 10432 8708 10434
rect 8477 10376 8482 10432
rect 8538 10376 8708 10432
rect 8477 10374 8708 10376
rect 8477 10371 8543 10374
rect 8702 10372 8708 10374
rect 8772 10372 8778 10436
rect 3165 10368 3481 10369
rect 0 10298 800 10328
rect 3165 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3481 10368
rect 3165 10303 3481 10304
rect 7604 10368 7920 10369
rect 7604 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7920 10368
rect 7604 10303 7920 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 7046 10236 7052 10300
rect 7116 10298 7122 10300
rect 7373 10298 7439 10301
rect 8848 10298 8908 10510
rect 10041 10507 10107 10510
rect 14038 10508 14044 10572
rect 14108 10570 14114 10572
rect 14733 10570 14799 10573
rect 16389 10570 16455 10573
rect 14108 10568 14799 10570
rect 14108 10512 14738 10568
rect 14794 10512 14799 10568
rect 14108 10510 14799 10512
rect 14108 10508 14114 10510
rect 14733 10507 14799 10510
rect 14920 10568 16455 10570
rect 14920 10512 16394 10568
rect 16450 10512 16455 10568
rect 14920 10510 16455 10512
rect 9438 10372 9444 10436
rect 9508 10434 9514 10436
rect 10961 10434 11027 10437
rect 9508 10432 11027 10434
rect 9508 10376 10966 10432
rect 11022 10376 11027 10432
rect 9508 10374 11027 10376
rect 9508 10372 9514 10374
rect 10961 10371 11027 10374
rect 12433 10434 12499 10437
rect 14457 10434 14523 10437
rect 12433 10432 14523 10434
rect 12433 10376 12438 10432
rect 12494 10376 14462 10432
rect 14518 10376 14523 10432
rect 12433 10374 14523 10376
rect 12433 10371 12499 10374
rect 14457 10371 14523 10374
rect 14641 10434 14707 10437
rect 14920 10434 14980 10510
rect 16389 10507 16455 10510
rect 14641 10432 14980 10434
rect 14641 10376 14646 10432
rect 14702 10376 14980 10432
rect 14641 10374 14980 10376
rect 14641 10371 14707 10374
rect 12043 10368 12359 10369
rect 12043 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12359 10368
rect 12043 10303 12359 10304
rect 16482 10368 16798 10369
rect 16482 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16798 10368
rect 16482 10303 16798 10304
rect 9305 10300 9371 10301
rect 7116 10296 7439 10298
rect 7116 10240 7378 10296
rect 7434 10240 7439 10296
rect 7116 10238 7439 10240
rect 7116 10236 7122 10238
rect 7373 10235 7439 10238
rect 8158 10238 8908 10298
rect 6637 10162 6703 10165
rect 8158 10162 8218 10238
rect 9254 10236 9260 10300
rect 9324 10298 9371 10300
rect 9765 10300 9831 10301
rect 9324 10296 9416 10298
rect 9366 10240 9416 10296
rect 9324 10238 9416 10240
rect 9765 10296 9812 10300
rect 9876 10298 9882 10300
rect 10317 10298 10383 10301
rect 11697 10298 11763 10301
rect 9765 10240 9770 10296
rect 9324 10236 9371 10238
rect 9305 10235 9371 10236
rect 9765 10236 9812 10240
rect 9876 10238 9922 10298
rect 10317 10296 11763 10298
rect 10317 10240 10322 10296
rect 10378 10240 11702 10296
rect 11758 10240 11763 10296
rect 10317 10238 11763 10240
rect 9876 10236 9882 10238
rect 9765 10235 9831 10236
rect 10317 10235 10383 10238
rect 11697 10235 11763 10238
rect 12433 10298 12499 10301
rect 14181 10298 14247 10301
rect 12433 10296 14247 10298
rect 12433 10240 12438 10296
rect 12494 10240 14186 10296
rect 14242 10240 14247 10296
rect 12433 10238 14247 10240
rect 12433 10235 12499 10238
rect 14181 10235 14247 10238
rect 6637 10160 8218 10162
rect 6637 10104 6642 10160
rect 6698 10104 8218 10160
rect 6637 10102 8218 10104
rect 8293 10162 8359 10165
rect 10777 10162 10843 10165
rect 11830 10162 11836 10164
rect 8293 10160 11836 10162
rect 8293 10104 8298 10160
rect 8354 10104 10782 10160
rect 10838 10104 11836 10160
rect 8293 10102 11836 10104
rect 6637 10099 6703 10102
rect 8293 10099 8359 10102
rect 10777 10099 10843 10102
rect 11830 10100 11836 10102
rect 11900 10162 11906 10164
rect 12801 10162 12867 10165
rect 11900 10160 12867 10162
rect 11900 10104 12806 10160
rect 12862 10104 12867 10160
rect 11900 10102 12867 10104
rect 11900 10100 11906 10102
rect 12801 10099 12867 10102
rect 12985 10162 13051 10165
rect 17585 10162 17651 10165
rect 12985 10160 17651 10162
rect 12985 10104 12990 10160
rect 13046 10104 17590 10160
rect 17646 10104 17651 10160
rect 12985 10102 17651 10104
rect 12985 10099 13051 10102
rect 17585 10099 17651 10102
rect 6913 10026 6979 10029
rect 7649 10026 7715 10029
rect 6913 10024 7715 10026
rect 6913 9968 6918 10024
rect 6974 9968 7654 10024
rect 7710 9968 7715 10024
rect 6913 9966 7715 9968
rect 6913 9963 6979 9966
rect 7649 9963 7715 9966
rect 8201 10026 8267 10029
rect 17033 10026 17099 10029
rect 8201 10024 17099 10026
rect 8201 9968 8206 10024
rect 8262 9968 17038 10024
rect 17094 9968 17099 10024
rect 8201 9966 17099 9968
rect 8201 9963 8267 9966
rect 17033 9963 17099 9966
rect 5441 9890 5507 9893
rect 7189 9890 7255 9893
rect 5441 9888 7255 9890
rect 5441 9832 5446 9888
rect 5502 9832 7194 9888
rect 7250 9832 7255 9888
rect 5441 9830 7255 9832
rect 5441 9827 5507 9830
rect 7189 9827 7255 9830
rect 8845 9890 8911 9893
rect 13445 9892 13511 9893
rect 8845 9888 12634 9890
rect 8845 9832 8850 9888
rect 8906 9832 12634 9888
rect 8845 9830 12634 9832
rect 8845 9827 8911 9830
rect 3825 9824 4141 9825
rect 3825 9760 3831 9824
rect 3895 9760 3911 9824
rect 3975 9760 3991 9824
rect 4055 9760 4071 9824
rect 4135 9760 4141 9824
rect 3825 9759 4141 9760
rect 8264 9824 8580 9825
rect 8264 9760 8270 9824
rect 8334 9760 8350 9824
rect 8414 9760 8430 9824
rect 8494 9760 8510 9824
rect 8574 9760 8580 9824
rect 8264 9759 8580 9760
rect 9806 9692 9812 9756
rect 9876 9754 9882 9756
rect 11513 9754 11579 9757
rect 9876 9752 11579 9754
rect 9876 9696 11518 9752
rect 11574 9696 11579 9752
rect 9876 9694 11579 9696
rect 9876 9692 9882 9694
rect 11513 9691 11579 9694
rect 0 9618 800 9648
rect 1945 9618 2011 9621
rect 0 9616 2011 9618
rect 0 9560 1950 9616
rect 2006 9560 2011 9616
rect 0 9558 2011 9560
rect 0 9528 800 9558
rect 1945 9555 2011 9558
rect 3417 9618 3483 9621
rect 3550 9618 3556 9620
rect 3417 9616 3556 9618
rect 3417 9560 3422 9616
rect 3478 9560 3556 9616
rect 3417 9558 3556 9560
rect 3417 9555 3483 9558
rect 3550 9556 3556 9558
rect 3620 9556 3626 9620
rect 4153 9618 4219 9621
rect 9121 9618 9187 9621
rect 4153 9616 9187 9618
rect 4153 9560 4158 9616
rect 4214 9560 9126 9616
rect 9182 9560 9187 9616
rect 4153 9558 9187 9560
rect 4153 9555 4219 9558
rect 9121 9555 9187 9558
rect 10225 9618 10291 9621
rect 11237 9618 11303 9621
rect 11697 9620 11763 9621
rect 11646 9618 11652 9620
rect 10225 9616 11303 9618
rect 10225 9560 10230 9616
rect 10286 9560 11242 9616
rect 11298 9560 11303 9616
rect 10225 9558 11303 9560
rect 11606 9558 11652 9618
rect 11716 9616 11763 9620
rect 11758 9560 11763 9616
rect 10225 9555 10291 9558
rect 11237 9555 11303 9558
rect 11646 9556 11652 9558
rect 11716 9556 11763 9560
rect 11697 9555 11763 9556
rect 11881 9618 11947 9621
rect 12433 9618 12499 9621
rect 11881 9616 12499 9618
rect 11881 9560 11886 9616
rect 11942 9560 12438 9616
rect 12494 9560 12499 9616
rect 11881 9558 12499 9560
rect 12574 9618 12634 9830
rect 13445 9888 13492 9892
rect 13556 9890 13562 9892
rect 13445 9832 13450 9888
rect 13445 9828 13492 9832
rect 13556 9830 13602 9890
rect 13556 9828 13562 9830
rect 13445 9827 13511 9828
rect 12703 9824 13019 9825
rect 12703 9760 12709 9824
rect 12773 9760 12789 9824
rect 12853 9760 12869 9824
rect 12933 9760 12949 9824
rect 13013 9760 13019 9824
rect 12703 9759 13019 9760
rect 17142 9824 17458 9825
rect 17142 9760 17148 9824
rect 17212 9760 17228 9824
rect 17292 9760 17308 9824
rect 17372 9760 17388 9824
rect 17452 9760 17458 9824
rect 17142 9759 17458 9760
rect 16941 9754 17007 9757
rect 13080 9752 17007 9754
rect 13080 9696 16946 9752
rect 17002 9696 17007 9752
rect 13080 9694 17007 9696
rect 13080 9618 13140 9694
rect 16941 9691 17007 9694
rect 14089 9620 14155 9621
rect 12574 9558 13140 9618
rect 11881 9555 11947 9558
rect 12433 9555 12499 9558
rect 14038 9556 14044 9620
rect 14108 9618 14155 9620
rect 16481 9618 16547 9621
rect 17769 9620 17835 9621
rect 17718 9618 17724 9620
rect 14108 9616 14200 9618
rect 14150 9560 14200 9616
rect 14108 9558 14200 9560
rect 14598 9616 16547 9618
rect 14598 9560 16486 9616
rect 16542 9560 16547 9616
rect 14598 9558 16547 9560
rect 17678 9558 17724 9618
rect 17788 9616 17835 9620
rect 17830 9560 17835 9616
rect 14108 9556 14155 9558
rect 14089 9555 14155 9556
rect 6177 9482 6243 9485
rect 6310 9482 6316 9484
rect 6177 9480 6316 9482
rect 6177 9424 6182 9480
rect 6238 9424 6316 9480
rect 6177 9422 6316 9424
rect 6177 9419 6243 9422
rect 6310 9420 6316 9422
rect 6380 9420 6386 9484
rect 6913 9482 6979 9485
rect 12985 9482 13051 9485
rect 6913 9480 13051 9482
rect 6913 9424 6918 9480
rect 6974 9424 12990 9480
rect 13046 9424 13051 9480
rect 6913 9422 13051 9424
rect 6913 9419 6979 9422
rect 12985 9419 13051 9422
rect 13997 9482 14063 9485
rect 14365 9482 14431 9485
rect 13997 9480 14431 9482
rect 13997 9424 14002 9480
rect 14058 9424 14370 9480
rect 14426 9424 14431 9480
rect 13997 9422 14431 9424
rect 13997 9419 14063 9422
rect 14365 9419 14431 9422
rect 12566 9284 12572 9348
rect 12636 9346 12642 9348
rect 13353 9346 13419 9349
rect 12636 9344 13419 9346
rect 12636 9288 13358 9344
rect 13414 9288 13419 9344
rect 12636 9286 13419 9288
rect 12636 9284 12642 9286
rect 13353 9283 13419 9286
rect 14365 9344 14431 9349
rect 14365 9288 14370 9344
rect 14426 9288 14431 9344
rect 14365 9283 14431 9288
rect 3165 9280 3481 9281
rect 3165 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3481 9280
rect 3165 9215 3481 9216
rect 7604 9280 7920 9281
rect 7604 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7920 9280
rect 7604 9215 7920 9216
rect 12043 9280 12359 9281
rect 12043 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12359 9280
rect 12043 9215 12359 9216
rect 4245 9210 4311 9213
rect 8385 9210 8451 9213
rect 10133 9210 10199 9213
rect 11237 9210 11303 9213
rect 4245 9208 4354 9210
rect 4245 9152 4250 9208
rect 4306 9152 4354 9208
rect 4245 9147 4354 9152
rect 8385 9208 10058 9210
rect 8385 9152 8390 9208
rect 8446 9152 10058 9208
rect 8385 9150 10058 9152
rect 8385 9147 8451 9150
rect 1485 9074 1551 9077
rect 1485 9072 1594 9074
rect 1485 9016 1490 9072
rect 1546 9016 1594 9072
rect 1485 9011 1594 9016
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 1534 8669 1594 9011
rect 4294 8941 4354 9147
rect 6494 9012 6500 9076
rect 6564 9074 6570 9076
rect 9581 9074 9647 9077
rect 6564 9072 9647 9074
rect 6564 9016 9586 9072
rect 9642 9016 9647 9072
rect 6564 9014 9647 9016
rect 9998 9074 10058 9150
rect 10133 9208 11303 9210
rect 10133 9152 10138 9208
rect 10194 9152 11242 9208
rect 11298 9152 11303 9208
rect 10133 9150 11303 9152
rect 10133 9147 10199 9150
rect 11237 9147 11303 9150
rect 11646 9148 11652 9212
rect 11716 9210 11722 9212
rect 11789 9210 11855 9213
rect 11716 9208 11855 9210
rect 11716 9152 11794 9208
rect 11850 9152 11855 9208
rect 11716 9150 11855 9152
rect 11716 9148 11722 9150
rect 11789 9147 11855 9150
rect 12617 9210 12683 9213
rect 14368 9210 14428 9283
rect 12617 9208 12956 9210
rect 12617 9152 12622 9208
rect 12678 9152 12956 9208
rect 12617 9150 12956 9152
rect 12617 9147 12683 9150
rect 12896 9108 12956 9150
rect 13080 9150 14428 9210
rect 13080 9108 13140 9150
rect 9998 9014 12818 9074
rect 12896 9048 13140 9108
rect 13813 9074 13879 9077
rect 14598 9074 14658 9558
rect 16481 9555 16547 9558
rect 17718 9556 17724 9558
rect 17788 9556 17835 9560
rect 17769 9555 17835 9556
rect 16021 9482 16087 9485
rect 16941 9482 17007 9485
rect 16021 9480 17007 9482
rect 16021 9424 16026 9480
rect 16082 9424 16946 9480
rect 17002 9424 17007 9480
rect 16021 9422 17007 9424
rect 16021 9419 16087 9422
rect 16941 9419 17007 9422
rect 16482 9280 16798 9281
rect 16482 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16798 9280
rect 16482 9215 16798 9216
rect 15193 9074 15259 9077
rect 18597 9074 18663 9077
rect 13813 9072 14658 9074
rect 6564 9012 6570 9014
rect 9581 9011 9647 9014
rect 4245 8936 4354 8941
rect 4245 8880 4250 8936
rect 4306 8880 4354 8936
rect 4245 8878 4354 8880
rect 4245 8875 4311 8878
rect 7230 8876 7236 8940
rect 7300 8938 7306 8940
rect 12758 8938 12818 9014
rect 13813 9016 13818 9072
rect 13874 9016 14658 9072
rect 13813 9014 14658 9016
rect 14736 9072 18663 9074
rect 14736 9016 15198 9072
rect 15254 9016 18602 9072
rect 18658 9016 18663 9072
rect 14736 9014 18663 9016
rect 13813 9011 13879 9014
rect 13445 8938 13511 8941
rect 14736 8938 14796 9014
rect 15193 9011 15259 9014
rect 18597 9011 18663 9014
rect 7300 8878 8770 8938
rect 12758 8878 13140 8938
rect 7300 8876 7306 8878
rect 5390 8740 5396 8804
rect 5460 8802 5466 8804
rect 7833 8802 7899 8805
rect 5460 8800 7899 8802
rect 5460 8744 7838 8800
rect 7894 8744 7899 8800
rect 5460 8742 7899 8744
rect 8710 8802 8770 8878
rect 11605 8802 11671 8805
rect 8710 8800 11671 8802
rect 8710 8744 11610 8800
rect 11666 8744 11671 8800
rect 8710 8742 11671 8744
rect 13080 8802 13140 8878
rect 13445 8936 14796 8938
rect 13445 8880 13450 8936
rect 13506 8880 14796 8936
rect 13445 8878 14796 8880
rect 15653 8938 15719 8941
rect 17309 8938 17375 8941
rect 15653 8936 17375 8938
rect 15653 8880 15658 8936
rect 15714 8880 17314 8936
rect 17370 8880 17375 8936
rect 15653 8878 17375 8880
rect 13445 8875 13511 8878
rect 15653 8875 15719 8878
rect 17309 8875 17375 8878
rect 13997 8802 14063 8805
rect 13080 8800 14063 8802
rect 13080 8744 14002 8800
rect 14058 8744 14063 8800
rect 13080 8742 14063 8744
rect 5460 8740 5466 8742
rect 7833 8739 7899 8742
rect 11605 8739 11671 8742
rect 13997 8739 14063 8742
rect 3825 8736 4141 8737
rect 3825 8672 3831 8736
rect 3895 8672 3911 8736
rect 3975 8672 3991 8736
rect 4055 8672 4071 8736
rect 4135 8672 4141 8736
rect 3825 8671 4141 8672
rect 8264 8736 8580 8737
rect 8264 8672 8270 8736
rect 8334 8672 8350 8736
rect 8414 8672 8430 8736
rect 8494 8672 8510 8736
rect 8574 8672 8580 8736
rect 8264 8671 8580 8672
rect 12703 8736 13019 8737
rect 12703 8672 12709 8736
rect 12773 8672 12789 8736
rect 12853 8672 12869 8736
rect 12933 8672 12949 8736
rect 13013 8672 13019 8736
rect 12703 8671 13019 8672
rect 17142 8736 17458 8737
rect 17142 8672 17148 8736
rect 17212 8672 17228 8736
rect 17292 8672 17308 8736
rect 17372 8672 17388 8736
rect 17452 8672 17458 8736
rect 17142 8671 17458 8672
rect 1485 8664 1594 8669
rect 1485 8608 1490 8664
rect 1546 8608 1594 8664
rect 1485 8606 1594 8608
rect 1485 8603 1551 8606
rect 6310 8604 6316 8668
rect 6380 8666 6386 8668
rect 7281 8666 7347 8669
rect 6380 8664 7347 8666
rect 6380 8608 7286 8664
rect 7342 8608 7347 8664
rect 6380 8606 7347 8608
rect 6380 8604 6386 8606
rect 7281 8603 7347 8606
rect 7414 8604 7420 8668
rect 7484 8666 7490 8668
rect 8109 8666 8175 8669
rect 7484 8664 8175 8666
rect 7484 8608 8114 8664
rect 8170 8608 8175 8664
rect 7484 8606 8175 8608
rect 7484 8604 7490 8606
rect 8109 8603 8175 8606
rect 11053 8666 11119 8669
rect 12525 8666 12591 8669
rect 11053 8664 12591 8666
rect 11053 8608 11058 8664
rect 11114 8608 12530 8664
rect 12586 8608 12591 8664
rect 11053 8606 12591 8608
rect 11053 8603 11119 8606
rect 12525 8603 12591 8606
rect 6913 8530 6979 8533
rect 19333 8530 19399 8533
rect 6913 8528 19399 8530
rect 6913 8472 6918 8528
rect 6974 8472 19338 8528
rect 19394 8472 19399 8528
rect 6913 8470 19399 8472
rect 6913 8467 6979 8470
rect 19333 8467 19399 8470
rect 2589 8394 2655 8397
rect 6913 8394 6979 8397
rect 7741 8394 7807 8397
rect 2589 8392 6979 8394
rect 2589 8336 2594 8392
rect 2650 8336 6918 8392
rect 6974 8336 6979 8392
rect 2589 8334 6979 8336
rect 2589 8331 2655 8334
rect 6913 8331 6979 8334
rect 7054 8392 7807 8394
rect 7054 8336 7746 8392
rect 7802 8336 7807 8392
rect 7054 8334 7807 8336
rect 0 8258 800 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 800 8198
rect 1577 8195 1643 8198
rect 4521 8258 4587 8261
rect 7054 8258 7114 8334
rect 7741 8331 7807 8334
rect 8109 8394 8175 8397
rect 9121 8394 9187 8397
rect 8109 8392 9187 8394
rect 8109 8336 8114 8392
rect 8170 8336 9126 8392
rect 9182 8336 9187 8392
rect 8109 8334 9187 8336
rect 8109 8331 8175 8334
rect 9121 8331 9187 8334
rect 11094 8332 11100 8396
rect 11164 8394 11170 8396
rect 13813 8394 13879 8397
rect 11164 8392 13879 8394
rect 11164 8336 13818 8392
rect 13874 8336 13879 8392
rect 11164 8334 13879 8336
rect 11164 8332 11170 8334
rect 13813 8331 13879 8334
rect 13997 8394 14063 8397
rect 14733 8394 14799 8397
rect 13997 8392 14799 8394
rect 13997 8336 14002 8392
rect 14058 8336 14738 8392
rect 14794 8336 14799 8392
rect 13997 8334 14799 8336
rect 13997 8331 14063 8334
rect 14733 8331 14799 8334
rect 16849 8394 16915 8397
rect 16982 8394 16988 8396
rect 16849 8392 16988 8394
rect 16849 8336 16854 8392
rect 16910 8336 16988 8392
rect 16849 8334 16988 8336
rect 16849 8331 16915 8334
rect 16982 8332 16988 8334
rect 17052 8332 17058 8396
rect 17493 8394 17559 8397
rect 18321 8394 18387 8397
rect 17493 8392 18387 8394
rect 17493 8336 17498 8392
rect 17554 8336 18326 8392
rect 18382 8336 18387 8392
rect 17493 8334 18387 8336
rect 17493 8331 17559 8334
rect 18321 8331 18387 8334
rect 4521 8256 7114 8258
rect 4521 8200 4526 8256
rect 4582 8200 7114 8256
rect 4521 8198 7114 8200
rect 9121 8258 9187 8261
rect 9990 8258 9996 8260
rect 9121 8256 9996 8258
rect 9121 8200 9126 8256
rect 9182 8200 9996 8256
rect 9121 8198 9996 8200
rect 4521 8195 4587 8198
rect 9121 8195 9187 8198
rect 9990 8196 9996 8198
rect 10060 8196 10066 8260
rect 12709 8258 12775 8261
rect 14038 8258 14044 8260
rect 12709 8256 14044 8258
rect 12709 8200 12714 8256
rect 12770 8200 14044 8256
rect 12709 8198 14044 8200
rect 12709 8195 12775 8198
rect 14038 8196 14044 8198
rect 14108 8196 14114 8260
rect 14774 8196 14780 8260
rect 14844 8258 14850 8260
rect 15009 8258 15075 8261
rect 14844 8256 15075 8258
rect 14844 8200 15014 8256
rect 15070 8200 15075 8256
rect 14844 8198 15075 8200
rect 14844 8196 14850 8198
rect 15009 8195 15075 8198
rect 3165 8192 3481 8193
rect 3165 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3481 8192
rect 3165 8127 3481 8128
rect 7604 8192 7920 8193
rect 7604 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7920 8192
rect 7604 8127 7920 8128
rect 12043 8192 12359 8193
rect 12043 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12359 8192
rect 12043 8127 12359 8128
rect 16482 8192 16798 8193
rect 16482 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16798 8192
rect 16482 8127 16798 8128
rect 4705 8122 4771 8125
rect 7097 8122 7163 8125
rect 4705 8120 7163 8122
rect 4705 8064 4710 8120
rect 4766 8064 7102 8120
rect 7158 8064 7163 8120
rect 4705 8062 7163 8064
rect 4705 8059 4771 8062
rect 7097 8059 7163 8062
rect 9397 8122 9463 8125
rect 11278 8122 11284 8124
rect 9397 8120 11284 8122
rect 9397 8064 9402 8120
rect 9458 8064 11284 8120
rect 9397 8062 11284 8064
rect 9397 8059 9463 8062
rect 11278 8060 11284 8062
rect 11348 8060 11354 8124
rect 12525 8122 12591 8125
rect 15561 8122 15627 8125
rect 12525 8120 15627 8122
rect 12525 8064 12530 8120
rect 12586 8064 15566 8120
rect 15622 8064 15627 8120
rect 12525 8062 15627 8064
rect 12525 8059 12591 8062
rect 15561 8059 15627 8062
rect 2681 7986 2747 7989
rect 3417 7986 3483 7989
rect 5625 7986 5691 7989
rect 2681 7984 5691 7986
rect 2681 7928 2686 7984
rect 2742 7928 3422 7984
rect 3478 7928 5630 7984
rect 5686 7928 5691 7984
rect 2681 7926 5691 7928
rect 2681 7923 2747 7926
rect 3417 7923 3483 7926
rect 5625 7923 5691 7926
rect 7097 7986 7163 7989
rect 12249 7986 12315 7989
rect 7097 7984 12315 7986
rect 7097 7928 7102 7984
rect 7158 7928 12254 7984
rect 12310 7928 12315 7984
rect 7097 7926 12315 7928
rect 7097 7923 7163 7926
rect 12249 7923 12315 7926
rect 12525 7986 12591 7989
rect 17033 7986 17099 7989
rect 12525 7984 17099 7986
rect 12525 7928 12530 7984
rect 12586 7928 17038 7984
rect 17094 7928 17099 7984
rect 12525 7926 17099 7928
rect 12525 7923 12591 7926
rect 17033 7923 17099 7926
rect 5165 7850 5231 7853
rect 12249 7850 12315 7853
rect 5165 7848 12315 7850
rect 5165 7792 5170 7848
rect 5226 7792 12254 7848
rect 12310 7792 12315 7848
rect 5165 7790 12315 7792
rect 5165 7787 5231 7790
rect 12249 7787 12315 7790
rect 12801 7850 12867 7853
rect 18045 7850 18111 7853
rect 12801 7848 18111 7850
rect 12801 7792 12806 7848
rect 12862 7792 18050 7848
rect 18106 7792 18111 7848
rect 12801 7790 18111 7792
rect 12801 7787 12867 7790
rect 18045 7787 18111 7790
rect 9029 7714 9095 7717
rect 12525 7714 12591 7717
rect 9029 7712 12591 7714
rect 9029 7656 9034 7712
rect 9090 7656 12530 7712
rect 12586 7656 12591 7712
rect 9029 7654 12591 7656
rect 9029 7651 9095 7654
rect 12525 7651 12591 7654
rect 13169 7714 13235 7717
rect 15101 7714 15167 7717
rect 16389 7714 16455 7717
rect 13169 7712 16455 7714
rect 13169 7656 13174 7712
rect 13230 7656 15106 7712
rect 15162 7656 16394 7712
rect 16450 7656 16455 7712
rect 13169 7654 16455 7656
rect 13169 7651 13235 7654
rect 15101 7651 15167 7654
rect 16389 7651 16455 7654
rect 3825 7648 4141 7649
rect 0 7578 800 7608
rect 3825 7584 3831 7648
rect 3895 7584 3911 7648
rect 3975 7584 3991 7648
rect 4055 7584 4071 7648
rect 4135 7584 4141 7648
rect 3825 7583 4141 7584
rect 8264 7648 8580 7649
rect 8264 7584 8270 7648
rect 8334 7584 8350 7648
rect 8414 7584 8430 7648
rect 8494 7584 8510 7648
rect 8574 7584 8580 7648
rect 8264 7583 8580 7584
rect 12703 7648 13019 7649
rect 12703 7584 12709 7648
rect 12773 7584 12789 7648
rect 12853 7584 12869 7648
rect 12933 7584 12949 7648
rect 13013 7584 13019 7648
rect 12703 7583 13019 7584
rect 17142 7648 17458 7649
rect 17142 7584 17148 7648
rect 17212 7584 17228 7648
rect 17292 7584 17308 7648
rect 17372 7584 17388 7648
rect 17452 7584 17458 7648
rect 17142 7583 17458 7584
rect 2129 7578 2195 7581
rect 0 7576 2195 7578
rect 0 7520 2134 7576
rect 2190 7520 2195 7576
rect 0 7518 2195 7520
rect 0 7488 800 7518
rect 2129 7515 2195 7518
rect 11513 7578 11579 7581
rect 11646 7578 11652 7580
rect 11513 7576 11652 7578
rect 11513 7520 11518 7576
rect 11574 7520 11652 7576
rect 11513 7518 11652 7520
rect 11513 7515 11579 7518
rect 11646 7516 11652 7518
rect 11716 7516 11722 7580
rect 11830 7516 11836 7580
rect 11900 7578 11906 7580
rect 12157 7578 12223 7581
rect 11900 7576 12223 7578
rect 11900 7520 12162 7576
rect 12218 7520 12223 7576
rect 11900 7518 12223 7520
rect 11900 7516 11906 7518
rect 12157 7515 12223 7518
rect 13486 7516 13492 7580
rect 13556 7578 13562 7580
rect 16389 7578 16455 7581
rect 13556 7576 16455 7578
rect 13556 7520 16394 7576
rect 16450 7520 16455 7576
rect 13556 7518 16455 7520
rect 13556 7516 13562 7518
rect 16389 7515 16455 7518
rect 1853 7442 1919 7445
rect 9029 7442 9095 7445
rect 17033 7442 17099 7445
rect 1853 7440 17099 7442
rect 1853 7384 1858 7440
rect 1914 7384 9034 7440
rect 9090 7384 17038 7440
rect 17094 7384 17099 7440
rect 1853 7382 17099 7384
rect 1853 7379 1919 7382
rect 9029 7379 9095 7382
rect 17033 7379 17099 7382
rect 2129 7306 2195 7309
rect 4613 7306 4679 7309
rect 13721 7306 13787 7309
rect 2129 7304 4679 7306
rect 2129 7248 2134 7304
rect 2190 7248 4618 7304
rect 4674 7248 4679 7304
rect 2129 7246 4679 7248
rect 2129 7243 2195 7246
rect 4613 7243 4679 7246
rect 7284 7304 13787 7306
rect 7284 7248 13726 7304
rect 13782 7248 13787 7304
rect 7284 7246 13787 7248
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 4337 7036 4403 7037
rect 4286 6972 4292 7036
rect 4356 7034 4403 7036
rect 4356 7032 4448 7034
rect 4398 6976 4448 7032
rect 4356 6974 4448 6976
rect 4356 6972 4403 6974
rect 4337 6971 4403 6972
rect 0 6898 800 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 800 6838
rect 1577 6835 1643 6838
rect 2405 6898 2471 6901
rect 5073 6898 5139 6901
rect 2405 6896 5139 6898
rect 2405 6840 2410 6896
rect 2466 6840 5078 6896
rect 5134 6840 5139 6896
rect 2405 6838 5139 6840
rect 2405 6835 2471 6838
rect 5073 6835 5139 6838
rect 6269 6898 6335 6901
rect 7284 6898 7344 7246
rect 13721 7243 13787 7246
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 13445 7034 13511 7037
rect 13670 7034 13676 7036
rect 13445 7032 13676 7034
rect 13445 6976 13450 7032
rect 13506 6976 13676 7032
rect 13445 6974 13676 6976
rect 13445 6971 13511 6974
rect 13670 6972 13676 6974
rect 13740 6972 13746 7036
rect 6269 6896 7344 6898
rect 6269 6840 6274 6896
rect 6330 6840 7344 6896
rect 6269 6838 7344 6840
rect 7465 6898 7531 6901
rect 12249 6898 12315 6901
rect 7465 6896 12315 6898
rect 7465 6840 7470 6896
rect 7526 6840 12254 6896
rect 12310 6840 12315 6896
rect 7465 6838 12315 6840
rect 6269 6835 6335 6838
rect 7465 6835 7531 6838
rect 12249 6835 12315 6838
rect 12433 6898 12499 6901
rect 13353 6898 13419 6901
rect 12433 6896 13419 6898
rect 12433 6840 12438 6896
rect 12494 6840 13358 6896
rect 13414 6840 13419 6896
rect 12433 6838 13419 6840
rect 12433 6835 12499 6838
rect 13353 6835 13419 6838
rect 14406 6836 14412 6900
rect 14476 6898 14482 6900
rect 14641 6898 14707 6901
rect 14476 6896 14707 6898
rect 14476 6840 14646 6896
rect 14702 6840 14707 6896
rect 14476 6838 14707 6840
rect 14476 6836 14482 6838
rect 14641 6835 14707 6838
rect 1342 6700 1348 6764
rect 1412 6762 1418 6764
rect 4061 6762 4127 6765
rect 1412 6760 4127 6762
rect 1412 6704 4066 6760
rect 4122 6704 4127 6760
rect 1412 6702 4127 6704
rect 1412 6700 1418 6702
rect 4061 6699 4127 6702
rect 5165 6762 5231 6765
rect 11094 6762 11100 6764
rect 5165 6760 11100 6762
rect 5165 6704 5170 6760
rect 5226 6704 11100 6760
rect 5165 6702 11100 6704
rect 5165 6699 5231 6702
rect 11094 6700 11100 6702
rect 11164 6700 11170 6764
rect 11462 6700 11468 6764
rect 11532 6762 11538 6764
rect 12617 6762 12683 6765
rect 11532 6760 12683 6762
rect 11532 6704 12622 6760
rect 12678 6704 12683 6760
rect 11532 6702 12683 6704
rect 11532 6700 11538 6702
rect 12617 6699 12683 6702
rect 7005 6626 7071 6629
rect 7649 6626 7715 6629
rect 7005 6624 7715 6626
rect 7005 6568 7010 6624
rect 7066 6568 7654 6624
rect 7710 6568 7715 6624
rect 7005 6566 7715 6568
rect 7005 6563 7071 6566
rect 7649 6563 7715 6566
rect 9857 6626 9923 6629
rect 12341 6626 12407 6629
rect 9857 6624 12407 6626
rect 9857 6568 9862 6624
rect 9918 6568 12346 6624
rect 12402 6568 12407 6624
rect 9857 6566 12407 6568
rect 9857 6563 9923 6566
rect 12341 6563 12407 6566
rect 3825 6560 4141 6561
rect 3825 6496 3831 6560
rect 3895 6496 3911 6560
rect 3975 6496 3991 6560
rect 4055 6496 4071 6560
rect 4135 6496 4141 6560
rect 3825 6495 4141 6496
rect 8264 6560 8580 6561
rect 8264 6496 8270 6560
rect 8334 6496 8350 6560
rect 8414 6496 8430 6560
rect 8494 6496 8510 6560
rect 8574 6496 8580 6560
rect 8264 6495 8580 6496
rect 12703 6560 13019 6561
rect 12703 6496 12709 6560
rect 12773 6496 12789 6560
rect 12853 6496 12869 6560
rect 12933 6496 12949 6560
rect 13013 6496 13019 6560
rect 12703 6495 13019 6496
rect 17142 6560 17458 6561
rect 17142 6496 17148 6560
rect 17212 6496 17228 6560
rect 17292 6496 17308 6560
rect 17372 6496 17388 6560
rect 17452 6496 17458 6560
rect 17142 6495 17458 6496
rect 5625 6490 5691 6493
rect 7005 6490 7071 6493
rect 9489 6492 9555 6493
rect 5625 6488 7071 6490
rect 5625 6432 5630 6488
rect 5686 6432 7010 6488
rect 7066 6432 7071 6488
rect 5625 6430 7071 6432
rect 5625 6427 5691 6430
rect 7005 6427 7071 6430
rect 9438 6428 9444 6492
rect 9508 6490 9555 6492
rect 9508 6488 9600 6490
rect 9550 6432 9600 6488
rect 9508 6430 9600 6432
rect 9508 6428 9555 6430
rect 11278 6428 11284 6492
rect 11348 6490 11354 6492
rect 12525 6490 12591 6493
rect 11348 6488 12591 6490
rect 11348 6432 12530 6488
rect 12586 6432 12591 6488
rect 11348 6430 12591 6432
rect 11348 6428 11354 6430
rect 9489 6427 9555 6428
rect 12525 6427 12591 6430
rect 2957 6354 3023 6357
rect 10174 6354 10180 6356
rect 2957 6352 10180 6354
rect 2957 6296 2962 6352
rect 3018 6296 10180 6352
rect 2957 6294 10180 6296
rect 2957 6291 3023 6294
rect 10174 6292 10180 6294
rect 10244 6292 10250 6356
rect 16941 6354 17007 6357
rect 17493 6356 17559 6357
rect 17493 6354 17540 6356
rect 10366 6352 17007 6354
rect 10366 6296 16946 6352
rect 17002 6296 17007 6352
rect 10366 6294 17007 6296
rect 17448 6352 17540 6354
rect 17448 6296 17498 6352
rect 17448 6294 17540 6296
rect 0 6218 800 6248
rect 2313 6218 2379 6221
rect 2589 6218 2655 6221
rect 3417 6218 3483 6221
rect 0 6128 858 6218
rect 2313 6216 3618 6218
rect 2313 6160 2318 6216
rect 2374 6160 2594 6216
rect 2650 6160 3422 6216
rect 3478 6160 3618 6216
rect 2313 6158 3618 6160
rect 2313 6155 2379 6158
rect 2589 6155 2655 6158
rect 3417 6155 3483 6158
rect 798 6085 858 6128
rect 798 6080 907 6085
rect 798 6024 846 6080
rect 902 6024 907 6080
rect 798 6022 907 6024
rect 3558 6082 3618 6158
rect 6678 6156 6684 6220
rect 6748 6218 6754 6220
rect 10366 6218 10426 6294
rect 16941 6291 17007 6294
rect 17493 6292 17540 6294
rect 17604 6292 17610 6356
rect 17493 6291 17559 6292
rect 6748 6158 10426 6218
rect 10961 6218 11027 6221
rect 14181 6218 14247 6221
rect 10961 6216 14247 6218
rect 10961 6160 10966 6216
rect 11022 6160 14186 6216
rect 14242 6160 14247 6216
rect 10961 6158 14247 6160
rect 6748 6156 6754 6158
rect 10961 6155 11027 6158
rect 14181 6155 14247 6158
rect 6913 6082 6979 6085
rect 12525 6084 12591 6085
rect 12525 6082 12572 6084
rect 3558 6080 6979 6082
rect 3558 6024 6918 6080
rect 6974 6024 6979 6080
rect 3558 6022 6979 6024
rect 12480 6080 12572 6082
rect 12480 6024 12530 6080
rect 12480 6022 12572 6024
rect 841 6019 907 6022
rect 6913 6019 6979 6022
rect 12525 6020 12572 6022
rect 12636 6020 12642 6084
rect 12801 6082 12867 6085
rect 13302 6082 13308 6084
rect 12801 6080 13308 6082
rect 12801 6024 12806 6080
rect 12862 6024 13308 6080
rect 12801 6022 13308 6024
rect 12525 6019 12591 6020
rect 12801 6019 12867 6022
rect 13302 6020 13308 6022
rect 13372 6020 13378 6084
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 8017 5946 8083 5949
rect 8477 5946 8543 5949
rect 8017 5944 8543 5946
rect 8017 5888 8022 5944
rect 8078 5888 8482 5944
rect 8538 5888 8543 5944
rect 8017 5886 8543 5888
rect 8017 5883 8083 5886
rect 8477 5883 8543 5886
rect 8661 5946 8727 5949
rect 8886 5946 8892 5948
rect 8661 5944 8892 5946
rect 8661 5888 8666 5944
rect 8722 5888 8892 5944
rect 8661 5886 8892 5888
rect 8661 5883 8727 5886
rect 8886 5884 8892 5886
rect 8956 5884 8962 5948
rect 13997 5946 14063 5949
rect 14590 5946 14596 5948
rect 13997 5944 14596 5946
rect 13997 5888 14002 5944
rect 14058 5888 14596 5944
rect 13997 5886 14596 5888
rect 13997 5883 14063 5886
rect 14590 5884 14596 5886
rect 14660 5884 14666 5948
rect 1669 5810 1735 5813
rect 9806 5810 9812 5812
rect 1669 5808 9812 5810
rect 1669 5752 1674 5808
rect 1730 5752 9812 5808
rect 1669 5750 9812 5752
rect 1669 5747 1735 5750
rect 9806 5748 9812 5750
rect 9876 5748 9882 5812
rect 10317 5810 10383 5813
rect 16389 5810 16455 5813
rect 10317 5808 16455 5810
rect 10317 5752 10322 5808
rect 10378 5752 16394 5808
rect 16450 5752 16455 5808
rect 10317 5750 16455 5752
rect 10317 5747 10383 5750
rect 16389 5747 16455 5750
rect 6269 5674 6335 5677
rect 6678 5674 6684 5676
rect 6269 5672 6684 5674
rect 6269 5616 6274 5672
rect 6330 5616 6684 5672
rect 6269 5614 6684 5616
rect 6269 5611 6335 5614
rect 6678 5612 6684 5614
rect 6748 5612 6754 5676
rect 8201 5674 8267 5677
rect 15469 5674 15535 5677
rect 16205 5674 16271 5677
rect 8201 5672 16271 5674
rect 8201 5616 8206 5672
rect 8262 5616 15474 5672
rect 15530 5616 16210 5672
rect 16266 5616 16271 5672
rect 8201 5614 16271 5616
rect 8201 5611 8267 5614
rect 15469 5611 15535 5614
rect 16205 5611 16271 5614
rect 0 5538 800 5568
rect 1577 5538 1643 5541
rect 0 5536 1643 5538
rect 0 5480 1582 5536
rect 1638 5480 1643 5536
rect 0 5478 1643 5480
rect 0 5448 800 5478
rect 1577 5475 1643 5478
rect 5390 5476 5396 5540
rect 5460 5538 5466 5540
rect 5533 5538 5599 5541
rect 10593 5540 10659 5541
rect 10542 5538 10548 5540
rect 5460 5536 5599 5538
rect 5460 5480 5538 5536
rect 5594 5480 5599 5536
rect 5460 5478 5599 5480
rect 10502 5478 10548 5538
rect 10612 5536 10659 5540
rect 10654 5480 10659 5536
rect 5460 5476 5466 5478
rect 5533 5475 5599 5478
rect 10542 5476 10548 5478
rect 10612 5476 10659 5480
rect 10593 5475 10659 5476
rect 3825 5472 4141 5473
rect 3825 5408 3831 5472
rect 3895 5408 3911 5472
rect 3975 5408 3991 5472
rect 4055 5408 4071 5472
rect 4135 5408 4141 5472
rect 3825 5407 4141 5408
rect 8264 5472 8580 5473
rect 8264 5408 8270 5472
rect 8334 5408 8350 5472
rect 8414 5408 8430 5472
rect 8494 5408 8510 5472
rect 8574 5408 8580 5472
rect 8264 5407 8580 5408
rect 12703 5472 13019 5473
rect 12703 5408 12709 5472
rect 12773 5408 12789 5472
rect 12853 5408 12869 5472
rect 12933 5408 12949 5472
rect 13013 5408 13019 5472
rect 12703 5407 13019 5408
rect 17142 5472 17458 5473
rect 17142 5408 17148 5472
rect 17212 5408 17228 5472
rect 17292 5408 17308 5472
rect 17372 5408 17388 5472
rect 17452 5408 17458 5472
rect 17142 5407 17458 5408
rect 2630 5204 2636 5268
rect 2700 5266 2706 5268
rect 3877 5266 3943 5269
rect 2700 5264 3943 5266
rect 2700 5208 3882 5264
rect 3938 5208 3943 5264
rect 2700 5206 3943 5208
rect 2700 5204 2706 5206
rect 3877 5203 3943 5206
rect 4153 5266 4219 5269
rect 6085 5266 6151 5269
rect 4153 5264 6151 5266
rect 4153 5208 4158 5264
rect 4214 5208 6090 5264
rect 6146 5208 6151 5264
rect 4153 5206 6151 5208
rect 4153 5203 4219 5206
rect 6085 5203 6151 5206
rect 7465 5266 7531 5269
rect 8702 5266 8708 5268
rect 7465 5264 8708 5266
rect 7465 5208 7470 5264
rect 7526 5208 8708 5264
rect 7465 5206 8708 5208
rect 7465 5203 7531 5206
rect 8702 5204 8708 5206
rect 8772 5204 8778 5268
rect 10041 5266 10107 5269
rect 16205 5266 16271 5269
rect 10041 5264 16271 5266
rect 10041 5208 10046 5264
rect 10102 5208 16210 5264
rect 16266 5208 16271 5264
rect 10041 5206 16271 5208
rect 10041 5203 10107 5206
rect 16205 5203 16271 5206
rect 2589 5130 2655 5133
rect 8017 5130 8083 5133
rect 17769 5130 17835 5133
rect 2589 5128 17835 5130
rect 2589 5072 2594 5128
rect 2650 5072 8022 5128
rect 8078 5072 17774 5128
rect 17830 5072 17835 5128
rect 2589 5070 17835 5072
rect 2589 5067 2655 5070
rect 8017 5067 8083 5070
rect 17769 5067 17835 5070
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 8017 4858 8083 4861
rect 8017 4856 10242 4858
rect 8017 4800 8022 4856
rect 8078 4800 10242 4856
rect 8017 4798 10242 4800
rect 0 4768 800 4798
rect 8017 4795 8083 4798
rect 1025 4722 1091 4725
rect 9397 4722 9463 4725
rect 1025 4720 9463 4722
rect 1025 4664 1030 4720
rect 1086 4664 9402 4720
rect 9458 4664 9463 4720
rect 1025 4662 9463 4664
rect 10182 4722 10242 4798
rect 16849 4722 16915 4725
rect 10182 4720 16915 4722
rect 10182 4664 16854 4720
rect 16910 4664 16915 4720
rect 10182 4662 16915 4664
rect 1025 4659 1091 4662
rect 9397 4659 9463 4662
rect 16849 4659 16915 4662
rect 4981 4588 5047 4589
rect 4981 4586 5028 4588
rect 4936 4584 5028 4586
rect 4936 4528 4986 4584
rect 4936 4526 5028 4528
rect 4981 4524 5028 4526
rect 5092 4524 5098 4588
rect 5165 4586 5231 4589
rect 5165 4584 12450 4586
rect 5165 4528 5170 4584
rect 5226 4528 12450 4584
rect 5165 4526 12450 4528
rect 4981 4523 5047 4524
rect 5165 4523 5231 4526
rect 6126 4388 6132 4452
rect 6196 4450 6202 4452
rect 8017 4450 8083 4453
rect 6196 4448 8083 4450
rect 6196 4392 8022 4448
rect 8078 4392 8083 4448
rect 6196 4390 8083 4392
rect 6196 4388 6202 4390
rect 8017 4387 8083 4390
rect 3825 4384 4141 4385
rect 3825 4320 3831 4384
rect 3895 4320 3911 4384
rect 3975 4320 3991 4384
rect 4055 4320 4071 4384
rect 4135 4320 4141 4384
rect 3825 4319 4141 4320
rect 8264 4384 8580 4385
rect 8264 4320 8270 4384
rect 8334 4320 8350 4384
rect 8414 4320 8430 4384
rect 8494 4320 8510 4384
rect 8574 4320 8580 4384
rect 8264 4319 8580 4320
rect 841 4314 907 4317
rect 798 4312 907 4314
rect 798 4256 846 4312
rect 902 4256 907 4312
rect 798 4251 907 4256
rect 798 4208 858 4251
rect 0 4118 858 4208
rect 2957 4180 3023 4181
rect 2957 4178 3004 4180
rect 2912 4176 3004 4178
rect 2912 4120 2962 4176
rect 2912 4118 3004 4120
rect 0 4088 800 4118
rect 2957 4116 3004 4118
rect 3068 4116 3074 4180
rect 9622 4116 9628 4180
rect 9692 4178 9698 4180
rect 10317 4178 10383 4181
rect 9692 4176 10383 4178
rect 9692 4120 10322 4176
rect 10378 4120 10383 4176
rect 9692 4118 10383 4120
rect 12390 4178 12450 4526
rect 12703 4384 13019 4385
rect 12703 4320 12709 4384
rect 12773 4320 12789 4384
rect 12853 4320 12869 4384
rect 12933 4320 12949 4384
rect 13013 4320 13019 4384
rect 12703 4319 13019 4320
rect 17142 4384 17458 4385
rect 17142 4320 17148 4384
rect 17212 4320 17228 4384
rect 17292 4320 17308 4384
rect 17372 4320 17388 4384
rect 17452 4320 17458 4384
rect 17142 4319 17458 4320
rect 12893 4178 12959 4181
rect 12390 4176 12959 4178
rect 12390 4120 12898 4176
rect 12954 4120 12959 4176
rect 12390 4118 12959 4120
rect 9692 4116 9698 4118
rect 2957 4115 3023 4116
rect 10317 4115 10383 4118
rect 12893 4115 12959 4118
rect 1158 3980 1164 4044
rect 1228 4042 1234 4044
rect 4429 4042 4495 4045
rect 1228 4040 4495 4042
rect 1228 3984 4434 4040
rect 4490 3984 4495 4040
rect 1228 3982 4495 3984
rect 1228 3980 1234 3982
rect 4429 3979 4495 3982
rect 8017 4042 8083 4045
rect 15377 4042 15443 4045
rect 8017 4040 15443 4042
rect 8017 3984 8022 4040
rect 8078 3984 15382 4040
rect 15438 3984 15443 4040
rect 8017 3982 15443 3984
rect 8017 3979 8083 3982
rect 15377 3979 15443 3982
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 6453 3772 6519 3773
rect 15469 3772 15535 3773
rect 790 3708 796 3772
rect 860 3770 866 3772
rect 6453 3770 6500 3772
rect 860 3710 2790 3770
rect 6408 3768 6500 3770
rect 6408 3712 6458 3768
rect 6408 3710 6500 3712
rect 860 3708 866 3710
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 2730 3634 2790 3710
rect 6453 3708 6500 3710
rect 6564 3708 6570 3772
rect 15469 3770 15516 3772
rect 15424 3768 15516 3770
rect 15424 3712 15474 3768
rect 15424 3710 15516 3712
rect 15469 3708 15516 3710
rect 15580 3708 15586 3772
rect 6453 3707 6519 3708
rect 15469 3707 15535 3708
rect 7833 3634 7899 3637
rect 2730 3632 7899 3634
rect 2730 3576 7838 3632
rect 7894 3576 7899 3632
rect 2730 3574 7899 3576
rect 7833 3571 7899 3574
rect 12341 3634 12407 3637
rect 14549 3634 14615 3637
rect 12341 3632 14615 3634
rect 12341 3576 12346 3632
rect 12402 3576 14554 3632
rect 14610 3576 14615 3632
rect 12341 3574 14615 3576
rect 12341 3571 12407 3574
rect 14549 3571 14615 3574
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 4429 3498 4495 3501
rect 5625 3498 5691 3501
rect 4429 3496 5691 3498
rect 4429 3440 4434 3496
rect 4490 3440 5630 3496
rect 5686 3440 5691 3496
rect 4429 3438 5691 3440
rect 0 3408 800 3438
rect 4429 3435 4495 3438
rect 5625 3435 5691 3438
rect 6085 3498 6151 3501
rect 15142 3498 15148 3500
rect 6085 3496 15148 3498
rect 6085 3440 6090 3496
rect 6146 3440 15148 3496
rect 6085 3438 15148 3440
rect 6085 3435 6151 3438
rect 15142 3436 15148 3438
rect 15212 3436 15218 3500
rect 3825 3296 4141 3297
rect 3825 3232 3831 3296
rect 3895 3232 3911 3296
rect 3975 3232 3991 3296
rect 4055 3232 4071 3296
rect 4135 3232 4141 3296
rect 3825 3231 4141 3232
rect 8264 3296 8580 3297
rect 8264 3232 8270 3296
rect 8334 3232 8350 3296
rect 8414 3232 8430 3296
rect 8494 3232 8510 3296
rect 8574 3232 8580 3296
rect 8264 3231 8580 3232
rect 12703 3296 13019 3297
rect 12703 3232 12709 3296
rect 12773 3232 12789 3296
rect 12853 3232 12869 3296
rect 12933 3232 12949 3296
rect 13013 3232 13019 3296
rect 12703 3231 13019 3232
rect 17142 3296 17458 3297
rect 17142 3232 17148 3296
rect 17212 3232 17228 3296
rect 17292 3232 17308 3296
rect 17372 3232 17388 3296
rect 17452 3232 17458 3296
rect 17142 3231 17458 3232
rect 17769 3226 17835 3229
rect 17902 3226 17908 3228
rect 17769 3224 17908 3226
rect 17769 3168 17774 3224
rect 17830 3168 17908 3224
rect 17769 3166 17908 3168
rect 17769 3163 17835 3166
rect 17902 3164 17908 3166
rect 17972 3164 17978 3228
rect 974 3028 980 3092
rect 1044 3090 1050 3092
rect 10685 3090 10751 3093
rect 1044 3088 10751 3090
rect 1044 3032 10690 3088
rect 10746 3032 10751 3088
rect 1044 3030 10751 3032
rect 1044 3028 1050 3030
rect 10685 3027 10751 3030
rect 11789 3090 11855 3093
rect 17309 3090 17375 3093
rect 11789 3088 17375 3090
rect 11789 3032 11794 3088
rect 11850 3032 17314 3088
rect 17370 3032 17375 3088
rect 11789 3030 17375 3032
rect 11789 3027 11855 3030
rect 17309 3027 17375 3030
rect 841 2954 907 2957
rect 798 2952 907 2954
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2891 907 2896
rect 11237 2954 11303 2957
rect 14958 2954 14964 2956
rect 11237 2952 14964 2954
rect 11237 2896 11242 2952
rect 11298 2896 14964 2952
rect 11237 2894 14964 2896
rect 11237 2891 11303 2894
rect 14958 2892 14964 2894
rect 15028 2892 15034 2956
rect 798 2848 858 2891
rect 0 2758 858 2848
rect 0 2728 800 2758
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 3825 2208 4141 2209
rect 0 2138 800 2168
rect 3825 2144 3831 2208
rect 3895 2144 3911 2208
rect 3975 2144 3991 2208
rect 4055 2144 4071 2208
rect 4135 2144 4141 2208
rect 3825 2143 4141 2144
rect 8264 2208 8580 2209
rect 8264 2144 8270 2208
rect 8334 2144 8350 2208
rect 8414 2144 8430 2208
rect 8494 2144 8510 2208
rect 8574 2144 8580 2208
rect 8264 2143 8580 2144
rect 12703 2208 13019 2209
rect 12703 2144 12709 2208
rect 12773 2144 12789 2208
rect 12853 2144 12869 2208
rect 12933 2144 12949 2208
rect 13013 2144 13019 2208
rect 12703 2143 13019 2144
rect 17142 2208 17458 2209
rect 17142 2144 17148 2208
rect 17212 2144 17228 2208
rect 17292 2144 17308 2208
rect 17372 2144 17388 2208
rect 17452 2144 17458 2208
rect 17142 2143 17458 2144
rect 2129 2138 2195 2141
rect 0 2136 2195 2138
rect 0 2080 2134 2136
rect 2190 2080 2195 2136
rect 0 2078 2195 2080
rect 0 2048 800 2078
rect 2129 2075 2195 2078
rect 841 1594 907 1597
rect 798 1592 907 1594
rect 798 1536 846 1592
rect 902 1536 907 1592
rect 798 1531 907 1536
rect 798 1488 858 1531
rect 0 1398 858 1488
rect 0 1368 800 1398
rect 0 778 800 808
rect 2773 778 2839 781
rect 0 776 2839 778
rect 0 720 2778 776
rect 2834 720 2839 776
rect 0 718 2839 720
rect 0 688 800 718
rect 2773 715 2839 718
rect 0 98 800 128
rect 2865 98 2931 101
rect 0 96 2931 98
rect 0 40 2870 96
rect 2926 40 2931 96
rect 0 38 2931 40
rect 0 8 800 38
rect 2865 35 2931 38
<< via3 >>
rect 9260 19756 9324 19820
rect 16988 18124 17052 18188
rect 1348 17988 1412 18052
rect 1164 17580 1228 17644
rect 3831 17436 3895 17440
rect 3831 17380 3835 17436
rect 3835 17380 3891 17436
rect 3891 17380 3895 17436
rect 3831 17376 3895 17380
rect 3911 17436 3975 17440
rect 3911 17380 3915 17436
rect 3915 17380 3971 17436
rect 3971 17380 3975 17436
rect 3911 17376 3975 17380
rect 3991 17436 4055 17440
rect 3991 17380 3995 17436
rect 3995 17380 4051 17436
rect 4051 17380 4055 17436
rect 3991 17376 4055 17380
rect 4071 17436 4135 17440
rect 4071 17380 4075 17436
rect 4075 17380 4131 17436
rect 4131 17380 4135 17436
rect 4071 17376 4135 17380
rect 8270 17436 8334 17440
rect 8270 17380 8274 17436
rect 8274 17380 8330 17436
rect 8330 17380 8334 17436
rect 8270 17376 8334 17380
rect 8350 17436 8414 17440
rect 8350 17380 8354 17436
rect 8354 17380 8410 17436
rect 8410 17380 8414 17436
rect 8350 17376 8414 17380
rect 8430 17436 8494 17440
rect 8430 17380 8434 17436
rect 8434 17380 8490 17436
rect 8490 17380 8494 17436
rect 8430 17376 8494 17380
rect 8510 17436 8574 17440
rect 8510 17380 8514 17436
rect 8514 17380 8570 17436
rect 8570 17380 8574 17436
rect 8510 17376 8574 17380
rect 12709 17436 12773 17440
rect 12709 17380 12713 17436
rect 12713 17380 12769 17436
rect 12769 17380 12773 17436
rect 12709 17376 12773 17380
rect 12789 17436 12853 17440
rect 12789 17380 12793 17436
rect 12793 17380 12849 17436
rect 12849 17380 12853 17436
rect 12789 17376 12853 17380
rect 12869 17436 12933 17440
rect 12869 17380 12873 17436
rect 12873 17380 12929 17436
rect 12929 17380 12933 17436
rect 12869 17376 12933 17380
rect 12949 17436 13013 17440
rect 12949 17380 12953 17436
rect 12953 17380 13009 17436
rect 13009 17380 13013 17436
rect 12949 17376 13013 17380
rect 17148 17436 17212 17440
rect 17148 17380 17152 17436
rect 17152 17380 17208 17436
rect 17208 17380 17212 17436
rect 17148 17376 17212 17380
rect 17228 17436 17292 17440
rect 17228 17380 17232 17436
rect 17232 17380 17288 17436
rect 17288 17380 17292 17436
rect 17228 17376 17292 17380
rect 17308 17436 17372 17440
rect 17308 17380 17312 17436
rect 17312 17380 17368 17436
rect 17368 17380 17372 17436
rect 17308 17376 17372 17380
rect 17388 17436 17452 17440
rect 17388 17380 17392 17436
rect 17392 17380 17448 17436
rect 17448 17380 17452 17436
rect 17388 17376 17452 17380
rect 17724 17036 17788 17100
rect 9076 16900 9140 16964
rect 3171 16892 3235 16896
rect 3171 16836 3175 16892
rect 3175 16836 3231 16892
rect 3231 16836 3235 16892
rect 3171 16832 3235 16836
rect 3251 16892 3315 16896
rect 3251 16836 3255 16892
rect 3255 16836 3311 16892
rect 3311 16836 3315 16892
rect 3251 16832 3315 16836
rect 3331 16892 3395 16896
rect 3331 16836 3335 16892
rect 3335 16836 3391 16892
rect 3391 16836 3395 16892
rect 3331 16832 3395 16836
rect 3411 16892 3475 16896
rect 3411 16836 3415 16892
rect 3415 16836 3471 16892
rect 3471 16836 3475 16892
rect 3411 16832 3475 16836
rect 7610 16892 7674 16896
rect 7610 16836 7614 16892
rect 7614 16836 7670 16892
rect 7670 16836 7674 16892
rect 7610 16832 7674 16836
rect 7690 16892 7754 16896
rect 7690 16836 7694 16892
rect 7694 16836 7750 16892
rect 7750 16836 7754 16892
rect 7690 16832 7754 16836
rect 7770 16892 7834 16896
rect 7770 16836 7774 16892
rect 7774 16836 7830 16892
rect 7830 16836 7834 16892
rect 7770 16832 7834 16836
rect 7850 16892 7914 16896
rect 7850 16836 7854 16892
rect 7854 16836 7910 16892
rect 7910 16836 7914 16892
rect 7850 16832 7914 16836
rect 12049 16892 12113 16896
rect 12049 16836 12053 16892
rect 12053 16836 12109 16892
rect 12109 16836 12113 16892
rect 12049 16832 12113 16836
rect 12129 16892 12193 16896
rect 12129 16836 12133 16892
rect 12133 16836 12189 16892
rect 12189 16836 12193 16892
rect 12129 16832 12193 16836
rect 12209 16892 12273 16896
rect 12209 16836 12213 16892
rect 12213 16836 12269 16892
rect 12269 16836 12273 16892
rect 12209 16832 12273 16836
rect 12289 16892 12353 16896
rect 12289 16836 12293 16892
rect 12293 16836 12349 16892
rect 12349 16836 12353 16892
rect 12289 16832 12353 16836
rect 16488 16892 16552 16896
rect 16488 16836 16492 16892
rect 16492 16836 16548 16892
rect 16548 16836 16552 16892
rect 16488 16832 16552 16836
rect 16568 16892 16632 16896
rect 16568 16836 16572 16892
rect 16572 16836 16628 16892
rect 16628 16836 16632 16892
rect 16568 16832 16632 16836
rect 16648 16892 16712 16896
rect 16648 16836 16652 16892
rect 16652 16836 16708 16892
rect 16708 16836 16712 16892
rect 16648 16832 16712 16836
rect 16728 16892 16792 16896
rect 16728 16836 16732 16892
rect 16732 16836 16788 16892
rect 16788 16836 16792 16892
rect 16728 16832 16792 16836
rect 3004 16628 3068 16692
rect 9628 16764 9692 16828
rect 2636 16492 2700 16556
rect 3831 16348 3895 16352
rect 3831 16292 3835 16348
rect 3835 16292 3891 16348
rect 3891 16292 3895 16348
rect 3831 16288 3895 16292
rect 3911 16348 3975 16352
rect 3911 16292 3915 16348
rect 3915 16292 3971 16348
rect 3971 16292 3975 16348
rect 3911 16288 3975 16292
rect 3991 16348 4055 16352
rect 3991 16292 3995 16348
rect 3995 16292 4051 16348
rect 4051 16292 4055 16348
rect 3991 16288 4055 16292
rect 4071 16348 4135 16352
rect 4071 16292 4075 16348
rect 4075 16292 4131 16348
rect 4131 16292 4135 16348
rect 4071 16288 4135 16292
rect 8270 16348 8334 16352
rect 8270 16292 8274 16348
rect 8274 16292 8330 16348
rect 8330 16292 8334 16348
rect 8270 16288 8334 16292
rect 8350 16348 8414 16352
rect 8350 16292 8354 16348
rect 8354 16292 8410 16348
rect 8410 16292 8414 16348
rect 8350 16288 8414 16292
rect 8430 16348 8494 16352
rect 8430 16292 8434 16348
rect 8434 16292 8490 16348
rect 8490 16292 8494 16348
rect 8430 16288 8494 16292
rect 8510 16348 8574 16352
rect 8510 16292 8514 16348
rect 8514 16292 8570 16348
rect 8570 16292 8574 16348
rect 8510 16288 8574 16292
rect 12709 16348 12773 16352
rect 12709 16292 12713 16348
rect 12713 16292 12769 16348
rect 12769 16292 12773 16348
rect 12709 16288 12773 16292
rect 12789 16348 12853 16352
rect 12789 16292 12793 16348
rect 12793 16292 12849 16348
rect 12849 16292 12853 16348
rect 12789 16288 12853 16292
rect 12869 16348 12933 16352
rect 12869 16292 12873 16348
rect 12873 16292 12929 16348
rect 12929 16292 12933 16348
rect 12869 16288 12933 16292
rect 12949 16348 13013 16352
rect 12949 16292 12953 16348
rect 12953 16292 13009 16348
rect 13009 16292 13013 16348
rect 12949 16288 13013 16292
rect 17148 16348 17212 16352
rect 17148 16292 17152 16348
rect 17152 16292 17208 16348
rect 17208 16292 17212 16348
rect 17148 16288 17212 16292
rect 17228 16348 17292 16352
rect 17228 16292 17232 16348
rect 17232 16292 17288 16348
rect 17288 16292 17292 16348
rect 17228 16288 17292 16292
rect 17308 16348 17372 16352
rect 17308 16292 17312 16348
rect 17312 16292 17368 16348
rect 17368 16292 17372 16348
rect 17308 16288 17372 16292
rect 17388 16348 17452 16352
rect 17388 16292 17392 16348
rect 17392 16292 17448 16348
rect 17448 16292 17452 16348
rect 17388 16288 17452 16292
rect 4476 16220 4540 16284
rect 9996 16220 10060 16284
rect 3556 16084 3620 16148
rect 14780 15948 14844 16012
rect 6868 15872 6932 15876
rect 6868 15816 6882 15872
rect 6882 15816 6932 15872
rect 6868 15812 6932 15816
rect 3171 15804 3235 15808
rect 3171 15748 3175 15804
rect 3175 15748 3231 15804
rect 3231 15748 3235 15804
rect 3171 15744 3235 15748
rect 3251 15804 3315 15808
rect 3251 15748 3255 15804
rect 3255 15748 3311 15804
rect 3311 15748 3315 15804
rect 3251 15744 3315 15748
rect 3331 15804 3395 15808
rect 3331 15748 3335 15804
rect 3335 15748 3391 15804
rect 3391 15748 3395 15804
rect 3331 15744 3395 15748
rect 3411 15804 3475 15808
rect 3411 15748 3415 15804
rect 3415 15748 3471 15804
rect 3471 15748 3475 15804
rect 3411 15744 3475 15748
rect 7610 15804 7674 15808
rect 7610 15748 7614 15804
rect 7614 15748 7670 15804
rect 7670 15748 7674 15804
rect 7610 15744 7674 15748
rect 7690 15804 7754 15808
rect 7690 15748 7694 15804
rect 7694 15748 7750 15804
rect 7750 15748 7754 15804
rect 7690 15744 7754 15748
rect 7770 15804 7834 15808
rect 7770 15748 7774 15804
rect 7774 15748 7830 15804
rect 7830 15748 7834 15804
rect 7770 15744 7834 15748
rect 7850 15804 7914 15808
rect 7850 15748 7854 15804
rect 7854 15748 7910 15804
rect 7910 15748 7914 15804
rect 7850 15744 7914 15748
rect 12049 15804 12113 15808
rect 12049 15748 12053 15804
rect 12053 15748 12109 15804
rect 12109 15748 12113 15804
rect 12049 15744 12113 15748
rect 12129 15804 12193 15808
rect 12129 15748 12133 15804
rect 12133 15748 12189 15804
rect 12189 15748 12193 15804
rect 12129 15744 12193 15748
rect 12209 15804 12273 15808
rect 12209 15748 12213 15804
rect 12213 15748 12269 15804
rect 12269 15748 12273 15804
rect 12209 15744 12273 15748
rect 12289 15804 12353 15808
rect 12289 15748 12293 15804
rect 12293 15748 12349 15804
rect 12349 15748 12353 15804
rect 12289 15744 12353 15748
rect 16488 15804 16552 15808
rect 16488 15748 16492 15804
rect 16492 15748 16548 15804
rect 16548 15748 16552 15804
rect 16488 15744 16552 15748
rect 16568 15804 16632 15808
rect 16568 15748 16572 15804
rect 16572 15748 16628 15804
rect 16628 15748 16632 15804
rect 16568 15744 16632 15748
rect 16648 15804 16712 15808
rect 16648 15748 16652 15804
rect 16652 15748 16708 15804
rect 16708 15748 16712 15804
rect 16648 15744 16712 15748
rect 16728 15804 16792 15808
rect 16728 15748 16732 15804
rect 16732 15748 16788 15804
rect 16788 15748 16792 15804
rect 16728 15744 16792 15748
rect 15516 15404 15580 15468
rect 14596 15328 14660 15332
rect 14596 15272 14610 15328
rect 14610 15272 14660 15328
rect 14596 15268 14660 15272
rect 3831 15260 3895 15264
rect 3831 15204 3835 15260
rect 3835 15204 3891 15260
rect 3891 15204 3895 15260
rect 3831 15200 3895 15204
rect 3911 15260 3975 15264
rect 3911 15204 3915 15260
rect 3915 15204 3971 15260
rect 3971 15204 3975 15260
rect 3911 15200 3975 15204
rect 3991 15260 4055 15264
rect 3991 15204 3995 15260
rect 3995 15204 4051 15260
rect 4051 15204 4055 15260
rect 3991 15200 4055 15204
rect 4071 15260 4135 15264
rect 4071 15204 4075 15260
rect 4075 15204 4131 15260
rect 4131 15204 4135 15260
rect 4071 15200 4135 15204
rect 8270 15260 8334 15264
rect 8270 15204 8274 15260
rect 8274 15204 8330 15260
rect 8330 15204 8334 15260
rect 8270 15200 8334 15204
rect 8350 15260 8414 15264
rect 8350 15204 8354 15260
rect 8354 15204 8410 15260
rect 8410 15204 8414 15260
rect 8350 15200 8414 15204
rect 8430 15260 8494 15264
rect 8430 15204 8434 15260
rect 8434 15204 8490 15260
rect 8490 15204 8494 15260
rect 8430 15200 8494 15204
rect 8510 15260 8574 15264
rect 8510 15204 8514 15260
rect 8514 15204 8570 15260
rect 8570 15204 8574 15260
rect 8510 15200 8574 15204
rect 12709 15260 12773 15264
rect 12709 15204 12713 15260
rect 12713 15204 12769 15260
rect 12769 15204 12773 15260
rect 12709 15200 12773 15204
rect 12789 15260 12853 15264
rect 12789 15204 12793 15260
rect 12793 15204 12849 15260
rect 12849 15204 12853 15260
rect 12789 15200 12853 15204
rect 12869 15260 12933 15264
rect 12869 15204 12873 15260
rect 12873 15204 12929 15260
rect 12929 15204 12933 15260
rect 12869 15200 12933 15204
rect 12949 15260 13013 15264
rect 12949 15204 12953 15260
rect 12953 15204 13009 15260
rect 13009 15204 13013 15260
rect 12949 15200 13013 15204
rect 17148 15260 17212 15264
rect 17148 15204 17152 15260
rect 17152 15204 17208 15260
rect 17208 15204 17212 15260
rect 17148 15200 17212 15204
rect 17228 15260 17292 15264
rect 17228 15204 17232 15260
rect 17232 15204 17288 15260
rect 17288 15204 17292 15260
rect 17228 15200 17292 15204
rect 17308 15260 17372 15264
rect 17308 15204 17312 15260
rect 17312 15204 17368 15260
rect 17368 15204 17372 15260
rect 17308 15200 17372 15204
rect 17388 15260 17452 15264
rect 17388 15204 17392 15260
rect 17392 15204 17448 15260
rect 17448 15204 17452 15260
rect 17388 15200 17452 15204
rect 7052 15132 7116 15196
rect 17908 14996 17972 15060
rect 8708 14724 8772 14788
rect 3171 14716 3235 14720
rect 3171 14660 3175 14716
rect 3175 14660 3231 14716
rect 3231 14660 3235 14716
rect 3171 14656 3235 14660
rect 3251 14716 3315 14720
rect 3251 14660 3255 14716
rect 3255 14660 3311 14716
rect 3311 14660 3315 14716
rect 3251 14656 3315 14660
rect 3331 14716 3395 14720
rect 3331 14660 3335 14716
rect 3335 14660 3391 14716
rect 3391 14660 3395 14716
rect 3331 14656 3395 14660
rect 3411 14716 3475 14720
rect 3411 14660 3415 14716
rect 3415 14660 3471 14716
rect 3471 14660 3475 14716
rect 3411 14656 3475 14660
rect 7610 14716 7674 14720
rect 7610 14660 7614 14716
rect 7614 14660 7670 14716
rect 7670 14660 7674 14716
rect 7610 14656 7674 14660
rect 7690 14716 7754 14720
rect 7690 14660 7694 14716
rect 7694 14660 7750 14716
rect 7750 14660 7754 14716
rect 7690 14656 7754 14660
rect 7770 14716 7834 14720
rect 7770 14660 7774 14716
rect 7774 14660 7830 14716
rect 7830 14660 7834 14716
rect 7770 14656 7834 14660
rect 7850 14716 7914 14720
rect 7850 14660 7854 14716
rect 7854 14660 7910 14716
rect 7910 14660 7914 14716
rect 7850 14656 7914 14660
rect 11468 14588 11532 14652
rect 11100 14452 11164 14516
rect 12049 14716 12113 14720
rect 12049 14660 12053 14716
rect 12053 14660 12109 14716
rect 12109 14660 12113 14716
rect 12049 14656 12113 14660
rect 12129 14716 12193 14720
rect 12129 14660 12133 14716
rect 12133 14660 12189 14716
rect 12189 14660 12193 14716
rect 12129 14656 12193 14660
rect 12209 14716 12273 14720
rect 12209 14660 12213 14716
rect 12213 14660 12269 14716
rect 12269 14660 12273 14716
rect 12209 14656 12273 14660
rect 12289 14716 12353 14720
rect 12289 14660 12293 14716
rect 12293 14660 12349 14716
rect 12349 14660 12353 14716
rect 12289 14656 12353 14660
rect 16488 14716 16552 14720
rect 16488 14660 16492 14716
rect 16492 14660 16548 14716
rect 16548 14660 16552 14716
rect 16488 14656 16552 14660
rect 16568 14716 16632 14720
rect 16568 14660 16572 14716
rect 16572 14660 16628 14716
rect 16628 14660 16632 14716
rect 16568 14656 16632 14660
rect 16648 14716 16712 14720
rect 16648 14660 16652 14716
rect 16652 14660 16708 14716
rect 16708 14660 16712 14716
rect 16648 14656 16712 14660
rect 16728 14716 16792 14720
rect 16728 14660 16732 14716
rect 16732 14660 16788 14716
rect 16788 14660 16792 14716
rect 16728 14656 16792 14660
rect 10732 14240 10796 14244
rect 10732 14184 10782 14240
rect 10782 14184 10796 14240
rect 10732 14180 10796 14184
rect 3831 14172 3895 14176
rect 3831 14116 3835 14172
rect 3835 14116 3891 14172
rect 3891 14116 3895 14172
rect 3831 14112 3895 14116
rect 3911 14172 3975 14176
rect 3911 14116 3915 14172
rect 3915 14116 3971 14172
rect 3971 14116 3975 14172
rect 3911 14112 3975 14116
rect 3991 14172 4055 14176
rect 3991 14116 3995 14172
rect 3995 14116 4051 14172
rect 4051 14116 4055 14172
rect 3991 14112 4055 14116
rect 4071 14172 4135 14176
rect 4071 14116 4075 14172
rect 4075 14116 4131 14172
rect 4131 14116 4135 14172
rect 4071 14112 4135 14116
rect 8270 14172 8334 14176
rect 8270 14116 8274 14172
rect 8274 14116 8330 14172
rect 8330 14116 8334 14172
rect 8270 14112 8334 14116
rect 8350 14172 8414 14176
rect 8350 14116 8354 14172
rect 8354 14116 8410 14172
rect 8410 14116 8414 14172
rect 8350 14112 8414 14116
rect 8430 14172 8494 14176
rect 8430 14116 8434 14172
rect 8434 14116 8490 14172
rect 8490 14116 8494 14172
rect 8430 14112 8494 14116
rect 8510 14172 8574 14176
rect 8510 14116 8514 14172
rect 8514 14116 8570 14172
rect 8570 14116 8574 14172
rect 8510 14112 8574 14116
rect 12709 14172 12773 14176
rect 12709 14116 12713 14172
rect 12713 14116 12769 14172
rect 12769 14116 12773 14172
rect 12709 14112 12773 14116
rect 12789 14172 12853 14176
rect 12789 14116 12793 14172
rect 12793 14116 12849 14172
rect 12849 14116 12853 14172
rect 12789 14112 12853 14116
rect 12869 14172 12933 14176
rect 12869 14116 12873 14172
rect 12873 14116 12929 14172
rect 12929 14116 12933 14172
rect 12869 14112 12933 14116
rect 12949 14172 13013 14176
rect 12949 14116 12953 14172
rect 12953 14116 13009 14172
rect 13009 14116 13013 14172
rect 12949 14112 13013 14116
rect 17148 14172 17212 14176
rect 17148 14116 17152 14172
rect 17152 14116 17208 14172
rect 17208 14116 17212 14172
rect 17148 14112 17212 14116
rect 17228 14172 17292 14176
rect 17228 14116 17232 14172
rect 17232 14116 17288 14172
rect 17288 14116 17292 14172
rect 17228 14112 17292 14116
rect 17308 14172 17372 14176
rect 17308 14116 17312 14172
rect 17312 14116 17368 14172
rect 17368 14116 17372 14172
rect 17308 14112 17372 14116
rect 17388 14172 17452 14176
rect 17388 14116 17392 14172
rect 17392 14116 17448 14172
rect 17448 14116 17452 14172
rect 17388 14112 17452 14116
rect 796 14044 860 14108
rect 4292 14104 4356 14108
rect 4292 14048 4342 14104
rect 4342 14048 4356 14104
rect 4292 14044 4356 14048
rect 4844 14044 4908 14108
rect 17540 14044 17604 14108
rect 10364 13908 10428 13972
rect 980 13772 1044 13836
rect 11836 13696 11900 13700
rect 13308 13772 13372 13836
rect 11836 13640 11850 13696
rect 11850 13640 11900 13696
rect 11836 13636 11900 13640
rect 14044 13636 14108 13700
rect 15148 13636 15212 13700
rect 3171 13628 3235 13632
rect 3171 13572 3175 13628
rect 3175 13572 3231 13628
rect 3231 13572 3235 13628
rect 3171 13568 3235 13572
rect 3251 13628 3315 13632
rect 3251 13572 3255 13628
rect 3255 13572 3311 13628
rect 3311 13572 3315 13628
rect 3251 13568 3315 13572
rect 3331 13628 3395 13632
rect 3331 13572 3335 13628
rect 3335 13572 3391 13628
rect 3391 13572 3395 13628
rect 3331 13568 3395 13572
rect 3411 13628 3475 13632
rect 3411 13572 3415 13628
rect 3415 13572 3471 13628
rect 3471 13572 3475 13628
rect 3411 13568 3475 13572
rect 7610 13628 7674 13632
rect 7610 13572 7614 13628
rect 7614 13572 7670 13628
rect 7670 13572 7674 13628
rect 7610 13568 7674 13572
rect 7690 13628 7754 13632
rect 7690 13572 7694 13628
rect 7694 13572 7750 13628
rect 7750 13572 7754 13628
rect 7690 13568 7754 13572
rect 7770 13628 7834 13632
rect 7770 13572 7774 13628
rect 7774 13572 7830 13628
rect 7830 13572 7834 13628
rect 7770 13568 7834 13572
rect 7850 13628 7914 13632
rect 7850 13572 7854 13628
rect 7854 13572 7910 13628
rect 7910 13572 7914 13628
rect 7850 13568 7914 13572
rect 12049 13628 12113 13632
rect 12049 13572 12053 13628
rect 12053 13572 12109 13628
rect 12109 13572 12113 13628
rect 12049 13568 12113 13572
rect 12129 13628 12193 13632
rect 12129 13572 12133 13628
rect 12133 13572 12189 13628
rect 12189 13572 12193 13628
rect 12129 13568 12193 13572
rect 12209 13628 12273 13632
rect 12209 13572 12213 13628
rect 12213 13572 12269 13628
rect 12269 13572 12273 13628
rect 12209 13568 12273 13572
rect 12289 13628 12353 13632
rect 12289 13572 12293 13628
rect 12293 13572 12349 13628
rect 12349 13572 12353 13628
rect 12289 13568 12353 13572
rect 16488 13628 16552 13632
rect 16488 13572 16492 13628
rect 16492 13572 16548 13628
rect 16548 13572 16552 13628
rect 16488 13568 16552 13572
rect 16568 13628 16632 13632
rect 16568 13572 16572 13628
rect 16572 13572 16628 13628
rect 16628 13572 16632 13628
rect 16568 13568 16632 13572
rect 16648 13628 16712 13632
rect 16648 13572 16652 13628
rect 16652 13572 16708 13628
rect 16708 13572 16712 13628
rect 16648 13568 16712 13572
rect 16728 13628 16792 13632
rect 16728 13572 16732 13628
rect 16732 13572 16788 13628
rect 16788 13572 16792 13628
rect 16728 13568 16792 13572
rect 6500 13500 6564 13564
rect 9444 13228 9508 13292
rect 7236 13092 7300 13156
rect 9812 13092 9876 13156
rect 3831 13084 3895 13088
rect 3831 13028 3835 13084
rect 3835 13028 3891 13084
rect 3891 13028 3895 13084
rect 3831 13024 3895 13028
rect 3911 13084 3975 13088
rect 3911 13028 3915 13084
rect 3915 13028 3971 13084
rect 3971 13028 3975 13084
rect 3911 13024 3975 13028
rect 3991 13084 4055 13088
rect 3991 13028 3995 13084
rect 3995 13028 4051 13084
rect 4051 13028 4055 13084
rect 3991 13024 4055 13028
rect 4071 13084 4135 13088
rect 4071 13028 4075 13084
rect 4075 13028 4131 13084
rect 4131 13028 4135 13084
rect 4071 13024 4135 13028
rect 8270 13084 8334 13088
rect 8270 13028 8274 13084
rect 8274 13028 8330 13084
rect 8330 13028 8334 13084
rect 8270 13024 8334 13028
rect 8350 13084 8414 13088
rect 8350 13028 8354 13084
rect 8354 13028 8410 13084
rect 8410 13028 8414 13084
rect 8350 13024 8414 13028
rect 8430 13084 8494 13088
rect 8430 13028 8434 13084
rect 8434 13028 8490 13084
rect 8490 13028 8494 13084
rect 8430 13024 8494 13028
rect 8510 13084 8574 13088
rect 8510 13028 8514 13084
rect 8514 13028 8570 13084
rect 8570 13028 8574 13084
rect 8510 13024 8574 13028
rect 12709 13084 12773 13088
rect 12709 13028 12713 13084
rect 12713 13028 12769 13084
rect 12769 13028 12773 13084
rect 12709 13024 12773 13028
rect 12789 13084 12853 13088
rect 12789 13028 12793 13084
rect 12793 13028 12849 13084
rect 12849 13028 12853 13084
rect 12789 13024 12853 13028
rect 12869 13084 12933 13088
rect 12869 13028 12873 13084
rect 12873 13028 12929 13084
rect 12929 13028 12933 13084
rect 12869 13024 12933 13028
rect 12949 13084 13013 13088
rect 12949 13028 12953 13084
rect 12953 13028 13009 13084
rect 13009 13028 13013 13084
rect 12949 13024 13013 13028
rect 17148 13084 17212 13088
rect 17148 13028 17152 13084
rect 17152 13028 17208 13084
rect 17208 13028 17212 13084
rect 17148 13024 17212 13028
rect 17228 13084 17292 13088
rect 17228 13028 17232 13084
rect 17232 13028 17288 13084
rect 17288 13028 17292 13084
rect 17228 13024 17292 13028
rect 17308 13084 17372 13088
rect 17308 13028 17312 13084
rect 17312 13028 17368 13084
rect 17368 13028 17372 13084
rect 17308 13024 17372 13028
rect 17388 13084 17452 13088
rect 17388 13028 17392 13084
rect 17392 13028 17448 13084
rect 17448 13028 17452 13084
rect 17388 13024 17452 13028
rect 3556 12684 3620 12748
rect 3171 12540 3235 12544
rect 3171 12484 3175 12540
rect 3175 12484 3231 12540
rect 3231 12484 3235 12540
rect 3171 12480 3235 12484
rect 3251 12540 3315 12544
rect 3251 12484 3255 12540
rect 3255 12484 3311 12540
rect 3311 12484 3315 12540
rect 3251 12480 3315 12484
rect 3331 12540 3395 12544
rect 3331 12484 3335 12540
rect 3335 12484 3391 12540
rect 3391 12484 3395 12540
rect 3331 12480 3395 12484
rect 3411 12540 3475 12544
rect 3411 12484 3415 12540
rect 3415 12484 3471 12540
rect 3471 12484 3475 12540
rect 3411 12480 3475 12484
rect 6132 12608 6196 12612
rect 6132 12552 6146 12608
rect 6146 12552 6196 12608
rect 6132 12548 6196 12552
rect 5028 12412 5092 12476
rect 7610 12540 7674 12544
rect 7610 12484 7614 12540
rect 7614 12484 7670 12540
rect 7670 12484 7674 12540
rect 7610 12480 7674 12484
rect 7690 12540 7754 12544
rect 7690 12484 7694 12540
rect 7694 12484 7750 12540
rect 7750 12484 7754 12540
rect 7690 12480 7754 12484
rect 7770 12540 7834 12544
rect 7770 12484 7774 12540
rect 7774 12484 7830 12540
rect 7830 12484 7834 12540
rect 7770 12480 7834 12484
rect 7850 12540 7914 12544
rect 7850 12484 7854 12540
rect 7854 12484 7910 12540
rect 7910 12484 7914 12540
rect 7850 12480 7914 12484
rect 9812 12548 9876 12612
rect 12049 12540 12113 12544
rect 12049 12484 12053 12540
rect 12053 12484 12109 12540
rect 12109 12484 12113 12540
rect 12049 12480 12113 12484
rect 12129 12540 12193 12544
rect 12129 12484 12133 12540
rect 12133 12484 12189 12540
rect 12189 12484 12193 12540
rect 12129 12480 12193 12484
rect 12209 12540 12273 12544
rect 12209 12484 12213 12540
rect 12213 12484 12269 12540
rect 12269 12484 12273 12540
rect 12209 12480 12273 12484
rect 12289 12540 12353 12544
rect 12289 12484 12293 12540
rect 12293 12484 12349 12540
rect 12349 12484 12353 12540
rect 12289 12480 12353 12484
rect 16488 12540 16552 12544
rect 16488 12484 16492 12540
rect 16492 12484 16548 12540
rect 16548 12484 16552 12540
rect 16488 12480 16552 12484
rect 16568 12540 16632 12544
rect 16568 12484 16572 12540
rect 16572 12484 16628 12540
rect 16628 12484 16632 12540
rect 16568 12480 16632 12484
rect 16648 12540 16712 12544
rect 16648 12484 16652 12540
rect 16652 12484 16708 12540
rect 16708 12484 16712 12540
rect 16648 12480 16712 12484
rect 16728 12540 16792 12544
rect 16728 12484 16732 12540
rect 16732 12484 16788 12540
rect 16788 12484 16792 12540
rect 16728 12480 16792 12484
rect 4292 12336 4356 12340
rect 4292 12280 4306 12336
rect 4306 12280 4356 12336
rect 4292 12276 4356 12280
rect 8708 12276 8772 12340
rect 9812 12276 9876 12340
rect 11652 12140 11716 12204
rect 6684 12004 6748 12068
rect 3831 11996 3895 12000
rect 3831 11940 3835 11996
rect 3835 11940 3891 11996
rect 3891 11940 3895 11996
rect 3831 11936 3895 11940
rect 3911 11996 3975 12000
rect 3911 11940 3915 11996
rect 3915 11940 3971 11996
rect 3971 11940 3975 11996
rect 3911 11936 3975 11940
rect 3991 11996 4055 12000
rect 3991 11940 3995 11996
rect 3995 11940 4051 11996
rect 4051 11940 4055 11996
rect 3991 11936 4055 11940
rect 4071 11996 4135 12000
rect 4071 11940 4075 11996
rect 4075 11940 4131 11996
rect 4131 11940 4135 11996
rect 4071 11936 4135 11940
rect 8270 11996 8334 12000
rect 8270 11940 8274 11996
rect 8274 11940 8330 11996
rect 8330 11940 8334 11996
rect 8270 11936 8334 11940
rect 8350 11996 8414 12000
rect 8350 11940 8354 11996
rect 8354 11940 8410 11996
rect 8410 11940 8414 11996
rect 8350 11936 8414 11940
rect 8430 11996 8494 12000
rect 8430 11940 8434 11996
rect 8434 11940 8490 11996
rect 8490 11940 8494 11996
rect 8430 11936 8494 11940
rect 8510 11996 8574 12000
rect 8510 11940 8514 11996
rect 8514 11940 8570 11996
rect 8570 11940 8574 11996
rect 8510 11936 8574 11940
rect 12709 11996 12773 12000
rect 12709 11940 12713 11996
rect 12713 11940 12769 11996
rect 12769 11940 12773 11996
rect 12709 11936 12773 11940
rect 12789 11996 12853 12000
rect 12789 11940 12793 11996
rect 12793 11940 12849 11996
rect 12849 11940 12853 11996
rect 12789 11936 12853 11940
rect 12869 11996 12933 12000
rect 12869 11940 12873 11996
rect 12873 11940 12929 11996
rect 12929 11940 12933 11996
rect 12869 11936 12933 11940
rect 12949 11996 13013 12000
rect 12949 11940 12953 11996
rect 12953 11940 13009 11996
rect 13009 11940 13013 11996
rect 12949 11936 13013 11940
rect 17148 11996 17212 12000
rect 17148 11940 17152 11996
rect 17152 11940 17208 11996
rect 17208 11940 17212 11996
rect 17148 11936 17212 11940
rect 17228 11996 17292 12000
rect 17228 11940 17232 11996
rect 17232 11940 17288 11996
rect 17288 11940 17292 11996
rect 17228 11936 17292 11940
rect 17308 11996 17372 12000
rect 17308 11940 17312 11996
rect 17312 11940 17368 11996
rect 17368 11940 17372 11996
rect 17308 11936 17372 11940
rect 17388 11996 17452 12000
rect 17388 11940 17392 11996
rect 17392 11940 17448 11996
rect 17448 11940 17452 11996
rect 17388 11936 17452 11940
rect 7420 11868 7484 11932
rect 9812 11868 9876 11932
rect 10180 11868 10244 11932
rect 13676 11868 13740 11932
rect 8892 11596 8956 11660
rect 10732 11460 10796 11524
rect 3171 11452 3235 11456
rect 3171 11396 3175 11452
rect 3175 11396 3231 11452
rect 3231 11396 3235 11452
rect 3171 11392 3235 11396
rect 3251 11452 3315 11456
rect 3251 11396 3255 11452
rect 3255 11396 3311 11452
rect 3311 11396 3315 11452
rect 3251 11392 3315 11396
rect 3331 11452 3395 11456
rect 3331 11396 3335 11452
rect 3335 11396 3391 11452
rect 3391 11396 3395 11452
rect 3331 11392 3395 11396
rect 3411 11452 3475 11456
rect 3411 11396 3415 11452
rect 3415 11396 3471 11452
rect 3471 11396 3475 11452
rect 3411 11392 3475 11396
rect 7610 11452 7674 11456
rect 7610 11396 7614 11452
rect 7614 11396 7670 11452
rect 7670 11396 7674 11452
rect 7610 11392 7674 11396
rect 7690 11452 7754 11456
rect 7690 11396 7694 11452
rect 7694 11396 7750 11452
rect 7750 11396 7754 11452
rect 7690 11392 7754 11396
rect 7770 11452 7834 11456
rect 7770 11396 7774 11452
rect 7774 11396 7830 11452
rect 7830 11396 7834 11452
rect 7770 11392 7834 11396
rect 7850 11452 7914 11456
rect 7850 11396 7854 11452
rect 7854 11396 7910 11452
rect 7910 11396 7914 11452
rect 7850 11392 7914 11396
rect 12049 11452 12113 11456
rect 12049 11396 12053 11452
rect 12053 11396 12109 11452
rect 12109 11396 12113 11452
rect 12049 11392 12113 11396
rect 12129 11452 12193 11456
rect 12129 11396 12133 11452
rect 12133 11396 12189 11452
rect 12189 11396 12193 11452
rect 12129 11392 12193 11396
rect 12209 11452 12273 11456
rect 12209 11396 12213 11452
rect 12213 11396 12269 11452
rect 12269 11396 12273 11452
rect 12209 11392 12273 11396
rect 12289 11452 12353 11456
rect 12289 11396 12293 11452
rect 12293 11396 12349 11452
rect 12349 11396 12353 11452
rect 12289 11392 12353 11396
rect 16488 11452 16552 11456
rect 16488 11396 16492 11452
rect 16492 11396 16548 11452
rect 16548 11396 16552 11452
rect 16488 11392 16552 11396
rect 16568 11452 16632 11456
rect 16568 11396 16572 11452
rect 16572 11396 16628 11452
rect 16628 11396 16632 11452
rect 16568 11392 16632 11396
rect 16648 11452 16712 11456
rect 16648 11396 16652 11452
rect 16652 11396 16708 11452
rect 16708 11396 16712 11452
rect 16648 11392 16712 11396
rect 16728 11452 16792 11456
rect 16728 11396 16732 11452
rect 16732 11396 16788 11452
rect 16788 11396 16792 11452
rect 16728 11392 16792 11396
rect 10548 11384 10612 11388
rect 10548 11328 10562 11384
rect 10562 11328 10612 11384
rect 10548 11324 10612 11328
rect 4844 11188 4908 11252
rect 8708 10916 8772 10980
rect 14412 11112 14476 11116
rect 14412 11056 14426 11112
rect 14426 11056 14476 11112
rect 14412 11052 14476 11056
rect 14964 11112 15028 11116
rect 14964 11056 14978 11112
rect 14978 11056 15028 11112
rect 14964 11052 15028 11056
rect 3831 10908 3895 10912
rect 3831 10852 3835 10908
rect 3835 10852 3891 10908
rect 3891 10852 3895 10908
rect 3831 10848 3895 10852
rect 3911 10908 3975 10912
rect 3911 10852 3915 10908
rect 3915 10852 3971 10908
rect 3971 10852 3975 10908
rect 3911 10848 3975 10852
rect 3991 10908 4055 10912
rect 3991 10852 3995 10908
rect 3995 10852 4051 10908
rect 4051 10852 4055 10908
rect 3991 10848 4055 10852
rect 4071 10908 4135 10912
rect 4071 10852 4075 10908
rect 4075 10852 4131 10908
rect 4131 10852 4135 10908
rect 4071 10848 4135 10852
rect 8270 10908 8334 10912
rect 8270 10852 8274 10908
rect 8274 10852 8330 10908
rect 8330 10852 8334 10908
rect 8270 10848 8334 10852
rect 8350 10908 8414 10912
rect 8350 10852 8354 10908
rect 8354 10852 8410 10908
rect 8410 10852 8414 10908
rect 8350 10848 8414 10852
rect 8430 10908 8494 10912
rect 8430 10852 8434 10908
rect 8434 10852 8490 10908
rect 8490 10852 8494 10908
rect 8430 10848 8494 10852
rect 8510 10908 8574 10912
rect 8510 10852 8514 10908
rect 8514 10852 8570 10908
rect 8570 10852 8574 10908
rect 8510 10848 8574 10852
rect 5396 10644 5460 10708
rect 4292 10508 4356 10572
rect 9076 10704 9140 10708
rect 9076 10648 9090 10704
rect 9090 10648 9140 10704
rect 9076 10644 9140 10648
rect 10364 10644 10428 10708
rect 11100 10644 11164 10708
rect 11836 10644 11900 10708
rect 12709 10908 12773 10912
rect 12709 10852 12713 10908
rect 12713 10852 12769 10908
rect 12769 10852 12773 10908
rect 12709 10848 12773 10852
rect 12789 10908 12853 10912
rect 12789 10852 12793 10908
rect 12793 10852 12849 10908
rect 12849 10852 12853 10908
rect 12789 10848 12853 10852
rect 12869 10908 12933 10912
rect 12869 10852 12873 10908
rect 12873 10852 12929 10908
rect 12929 10852 12933 10908
rect 12869 10848 12933 10852
rect 12949 10908 13013 10912
rect 12949 10852 12953 10908
rect 12953 10852 13009 10908
rect 13009 10852 13013 10908
rect 12949 10848 13013 10852
rect 17148 10908 17212 10912
rect 17148 10852 17152 10908
rect 17152 10852 17208 10908
rect 17208 10852 17212 10908
rect 17148 10848 17212 10852
rect 17228 10908 17292 10912
rect 17228 10852 17232 10908
rect 17232 10852 17288 10908
rect 17288 10852 17292 10908
rect 17228 10848 17292 10852
rect 17308 10908 17372 10912
rect 17308 10852 17312 10908
rect 17312 10852 17368 10908
rect 17368 10852 17372 10908
rect 17308 10848 17372 10852
rect 17388 10908 17452 10912
rect 17388 10852 17392 10908
rect 17392 10852 17448 10908
rect 17448 10852 17452 10908
rect 17388 10848 17452 10852
rect 4476 10372 4540 10436
rect 6868 10372 6932 10436
rect 8708 10372 8772 10436
rect 3171 10364 3235 10368
rect 3171 10308 3175 10364
rect 3175 10308 3231 10364
rect 3231 10308 3235 10364
rect 3171 10304 3235 10308
rect 3251 10364 3315 10368
rect 3251 10308 3255 10364
rect 3255 10308 3311 10364
rect 3311 10308 3315 10364
rect 3251 10304 3315 10308
rect 3331 10364 3395 10368
rect 3331 10308 3335 10364
rect 3335 10308 3391 10364
rect 3391 10308 3395 10364
rect 3331 10304 3395 10308
rect 3411 10364 3475 10368
rect 3411 10308 3415 10364
rect 3415 10308 3471 10364
rect 3471 10308 3475 10364
rect 3411 10304 3475 10308
rect 7610 10364 7674 10368
rect 7610 10308 7614 10364
rect 7614 10308 7670 10364
rect 7670 10308 7674 10364
rect 7610 10304 7674 10308
rect 7690 10364 7754 10368
rect 7690 10308 7694 10364
rect 7694 10308 7750 10364
rect 7750 10308 7754 10364
rect 7690 10304 7754 10308
rect 7770 10364 7834 10368
rect 7770 10308 7774 10364
rect 7774 10308 7830 10364
rect 7830 10308 7834 10364
rect 7770 10304 7834 10308
rect 7850 10364 7914 10368
rect 7850 10308 7854 10364
rect 7854 10308 7910 10364
rect 7910 10308 7914 10364
rect 7850 10304 7914 10308
rect 7052 10236 7116 10300
rect 14044 10508 14108 10572
rect 9444 10372 9508 10436
rect 12049 10364 12113 10368
rect 12049 10308 12053 10364
rect 12053 10308 12109 10364
rect 12109 10308 12113 10364
rect 12049 10304 12113 10308
rect 12129 10364 12193 10368
rect 12129 10308 12133 10364
rect 12133 10308 12189 10364
rect 12189 10308 12193 10364
rect 12129 10304 12193 10308
rect 12209 10364 12273 10368
rect 12209 10308 12213 10364
rect 12213 10308 12269 10364
rect 12269 10308 12273 10364
rect 12209 10304 12273 10308
rect 12289 10364 12353 10368
rect 12289 10308 12293 10364
rect 12293 10308 12349 10364
rect 12349 10308 12353 10364
rect 12289 10304 12353 10308
rect 16488 10364 16552 10368
rect 16488 10308 16492 10364
rect 16492 10308 16548 10364
rect 16548 10308 16552 10364
rect 16488 10304 16552 10308
rect 16568 10364 16632 10368
rect 16568 10308 16572 10364
rect 16572 10308 16628 10364
rect 16628 10308 16632 10364
rect 16568 10304 16632 10308
rect 16648 10364 16712 10368
rect 16648 10308 16652 10364
rect 16652 10308 16708 10364
rect 16708 10308 16712 10364
rect 16648 10304 16712 10308
rect 16728 10364 16792 10368
rect 16728 10308 16732 10364
rect 16732 10308 16788 10364
rect 16788 10308 16792 10364
rect 16728 10304 16792 10308
rect 9260 10296 9324 10300
rect 9260 10240 9310 10296
rect 9310 10240 9324 10296
rect 9260 10236 9324 10240
rect 9812 10296 9876 10300
rect 9812 10240 9826 10296
rect 9826 10240 9876 10296
rect 9812 10236 9876 10240
rect 11836 10100 11900 10164
rect 3831 9820 3895 9824
rect 3831 9764 3835 9820
rect 3835 9764 3891 9820
rect 3891 9764 3895 9820
rect 3831 9760 3895 9764
rect 3911 9820 3975 9824
rect 3911 9764 3915 9820
rect 3915 9764 3971 9820
rect 3971 9764 3975 9820
rect 3911 9760 3975 9764
rect 3991 9820 4055 9824
rect 3991 9764 3995 9820
rect 3995 9764 4051 9820
rect 4051 9764 4055 9820
rect 3991 9760 4055 9764
rect 4071 9820 4135 9824
rect 4071 9764 4075 9820
rect 4075 9764 4131 9820
rect 4131 9764 4135 9820
rect 4071 9760 4135 9764
rect 8270 9820 8334 9824
rect 8270 9764 8274 9820
rect 8274 9764 8330 9820
rect 8330 9764 8334 9820
rect 8270 9760 8334 9764
rect 8350 9820 8414 9824
rect 8350 9764 8354 9820
rect 8354 9764 8410 9820
rect 8410 9764 8414 9820
rect 8350 9760 8414 9764
rect 8430 9820 8494 9824
rect 8430 9764 8434 9820
rect 8434 9764 8490 9820
rect 8490 9764 8494 9820
rect 8430 9760 8494 9764
rect 8510 9820 8574 9824
rect 8510 9764 8514 9820
rect 8514 9764 8570 9820
rect 8570 9764 8574 9820
rect 8510 9760 8574 9764
rect 9812 9692 9876 9756
rect 3556 9556 3620 9620
rect 11652 9616 11716 9620
rect 11652 9560 11702 9616
rect 11702 9560 11716 9616
rect 11652 9556 11716 9560
rect 13492 9888 13556 9892
rect 13492 9832 13506 9888
rect 13506 9832 13556 9888
rect 13492 9828 13556 9832
rect 12709 9820 12773 9824
rect 12709 9764 12713 9820
rect 12713 9764 12769 9820
rect 12769 9764 12773 9820
rect 12709 9760 12773 9764
rect 12789 9820 12853 9824
rect 12789 9764 12793 9820
rect 12793 9764 12849 9820
rect 12849 9764 12853 9820
rect 12789 9760 12853 9764
rect 12869 9820 12933 9824
rect 12869 9764 12873 9820
rect 12873 9764 12929 9820
rect 12929 9764 12933 9820
rect 12869 9760 12933 9764
rect 12949 9820 13013 9824
rect 12949 9764 12953 9820
rect 12953 9764 13009 9820
rect 13009 9764 13013 9820
rect 12949 9760 13013 9764
rect 17148 9820 17212 9824
rect 17148 9764 17152 9820
rect 17152 9764 17208 9820
rect 17208 9764 17212 9820
rect 17148 9760 17212 9764
rect 17228 9820 17292 9824
rect 17228 9764 17232 9820
rect 17232 9764 17288 9820
rect 17288 9764 17292 9820
rect 17228 9760 17292 9764
rect 17308 9820 17372 9824
rect 17308 9764 17312 9820
rect 17312 9764 17368 9820
rect 17368 9764 17372 9820
rect 17308 9760 17372 9764
rect 17388 9820 17452 9824
rect 17388 9764 17392 9820
rect 17392 9764 17448 9820
rect 17448 9764 17452 9820
rect 17388 9760 17452 9764
rect 14044 9616 14108 9620
rect 14044 9560 14094 9616
rect 14094 9560 14108 9616
rect 14044 9556 14108 9560
rect 17724 9616 17788 9620
rect 17724 9560 17774 9616
rect 17774 9560 17788 9616
rect 6316 9420 6380 9484
rect 12572 9284 12636 9348
rect 3171 9276 3235 9280
rect 3171 9220 3175 9276
rect 3175 9220 3231 9276
rect 3231 9220 3235 9276
rect 3171 9216 3235 9220
rect 3251 9276 3315 9280
rect 3251 9220 3255 9276
rect 3255 9220 3311 9276
rect 3311 9220 3315 9276
rect 3251 9216 3315 9220
rect 3331 9276 3395 9280
rect 3331 9220 3335 9276
rect 3335 9220 3391 9276
rect 3391 9220 3395 9276
rect 3331 9216 3395 9220
rect 3411 9276 3475 9280
rect 3411 9220 3415 9276
rect 3415 9220 3471 9276
rect 3471 9220 3475 9276
rect 3411 9216 3475 9220
rect 7610 9276 7674 9280
rect 7610 9220 7614 9276
rect 7614 9220 7670 9276
rect 7670 9220 7674 9276
rect 7610 9216 7674 9220
rect 7690 9276 7754 9280
rect 7690 9220 7694 9276
rect 7694 9220 7750 9276
rect 7750 9220 7754 9276
rect 7690 9216 7754 9220
rect 7770 9276 7834 9280
rect 7770 9220 7774 9276
rect 7774 9220 7830 9276
rect 7830 9220 7834 9276
rect 7770 9216 7834 9220
rect 7850 9276 7914 9280
rect 7850 9220 7854 9276
rect 7854 9220 7910 9276
rect 7910 9220 7914 9276
rect 7850 9216 7914 9220
rect 12049 9276 12113 9280
rect 12049 9220 12053 9276
rect 12053 9220 12109 9276
rect 12109 9220 12113 9276
rect 12049 9216 12113 9220
rect 12129 9276 12193 9280
rect 12129 9220 12133 9276
rect 12133 9220 12189 9276
rect 12189 9220 12193 9276
rect 12129 9216 12193 9220
rect 12209 9276 12273 9280
rect 12209 9220 12213 9276
rect 12213 9220 12269 9276
rect 12269 9220 12273 9276
rect 12209 9216 12273 9220
rect 12289 9276 12353 9280
rect 12289 9220 12293 9276
rect 12293 9220 12349 9276
rect 12349 9220 12353 9276
rect 12289 9216 12353 9220
rect 6500 9012 6564 9076
rect 11652 9148 11716 9212
rect 17724 9556 17788 9560
rect 16488 9276 16552 9280
rect 16488 9220 16492 9276
rect 16492 9220 16548 9276
rect 16548 9220 16552 9276
rect 16488 9216 16552 9220
rect 16568 9276 16632 9280
rect 16568 9220 16572 9276
rect 16572 9220 16628 9276
rect 16628 9220 16632 9276
rect 16568 9216 16632 9220
rect 16648 9276 16712 9280
rect 16648 9220 16652 9276
rect 16652 9220 16708 9276
rect 16708 9220 16712 9276
rect 16648 9216 16712 9220
rect 16728 9276 16792 9280
rect 16728 9220 16732 9276
rect 16732 9220 16788 9276
rect 16788 9220 16792 9276
rect 16728 9216 16792 9220
rect 7236 8876 7300 8940
rect 5396 8740 5460 8804
rect 3831 8732 3895 8736
rect 3831 8676 3835 8732
rect 3835 8676 3891 8732
rect 3891 8676 3895 8732
rect 3831 8672 3895 8676
rect 3911 8732 3975 8736
rect 3911 8676 3915 8732
rect 3915 8676 3971 8732
rect 3971 8676 3975 8732
rect 3911 8672 3975 8676
rect 3991 8732 4055 8736
rect 3991 8676 3995 8732
rect 3995 8676 4051 8732
rect 4051 8676 4055 8732
rect 3991 8672 4055 8676
rect 4071 8732 4135 8736
rect 4071 8676 4075 8732
rect 4075 8676 4131 8732
rect 4131 8676 4135 8732
rect 4071 8672 4135 8676
rect 8270 8732 8334 8736
rect 8270 8676 8274 8732
rect 8274 8676 8330 8732
rect 8330 8676 8334 8732
rect 8270 8672 8334 8676
rect 8350 8732 8414 8736
rect 8350 8676 8354 8732
rect 8354 8676 8410 8732
rect 8410 8676 8414 8732
rect 8350 8672 8414 8676
rect 8430 8732 8494 8736
rect 8430 8676 8434 8732
rect 8434 8676 8490 8732
rect 8490 8676 8494 8732
rect 8430 8672 8494 8676
rect 8510 8732 8574 8736
rect 8510 8676 8514 8732
rect 8514 8676 8570 8732
rect 8570 8676 8574 8732
rect 8510 8672 8574 8676
rect 12709 8732 12773 8736
rect 12709 8676 12713 8732
rect 12713 8676 12769 8732
rect 12769 8676 12773 8732
rect 12709 8672 12773 8676
rect 12789 8732 12853 8736
rect 12789 8676 12793 8732
rect 12793 8676 12849 8732
rect 12849 8676 12853 8732
rect 12789 8672 12853 8676
rect 12869 8732 12933 8736
rect 12869 8676 12873 8732
rect 12873 8676 12929 8732
rect 12929 8676 12933 8732
rect 12869 8672 12933 8676
rect 12949 8732 13013 8736
rect 12949 8676 12953 8732
rect 12953 8676 13009 8732
rect 13009 8676 13013 8732
rect 12949 8672 13013 8676
rect 17148 8732 17212 8736
rect 17148 8676 17152 8732
rect 17152 8676 17208 8732
rect 17208 8676 17212 8732
rect 17148 8672 17212 8676
rect 17228 8732 17292 8736
rect 17228 8676 17232 8732
rect 17232 8676 17288 8732
rect 17288 8676 17292 8732
rect 17228 8672 17292 8676
rect 17308 8732 17372 8736
rect 17308 8676 17312 8732
rect 17312 8676 17368 8732
rect 17368 8676 17372 8732
rect 17308 8672 17372 8676
rect 17388 8732 17452 8736
rect 17388 8676 17392 8732
rect 17392 8676 17448 8732
rect 17448 8676 17452 8732
rect 17388 8672 17452 8676
rect 6316 8604 6380 8668
rect 7420 8604 7484 8668
rect 11100 8332 11164 8396
rect 16988 8332 17052 8396
rect 9996 8196 10060 8260
rect 14044 8196 14108 8260
rect 14780 8196 14844 8260
rect 3171 8188 3235 8192
rect 3171 8132 3175 8188
rect 3175 8132 3231 8188
rect 3231 8132 3235 8188
rect 3171 8128 3235 8132
rect 3251 8188 3315 8192
rect 3251 8132 3255 8188
rect 3255 8132 3311 8188
rect 3311 8132 3315 8188
rect 3251 8128 3315 8132
rect 3331 8188 3395 8192
rect 3331 8132 3335 8188
rect 3335 8132 3391 8188
rect 3391 8132 3395 8188
rect 3331 8128 3395 8132
rect 3411 8188 3475 8192
rect 3411 8132 3415 8188
rect 3415 8132 3471 8188
rect 3471 8132 3475 8188
rect 3411 8128 3475 8132
rect 7610 8188 7674 8192
rect 7610 8132 7614 8188
rect 7614 8132 7670 8188
rect 7670 8132 7674 8188
rect 7610 8128 7674 8132
rect 7690 8188 7754 8192
rect 7690 8132 7694 8188
rect 7694 8132 7750 8188
rect 7750 8132 7754 8188
rect 7690 8128 7754 8132
rect 7770 8188 7834 8192
rect 7770 8132 7774 8188
rect 7774 8132 7830 8188
rect 7830 8132 7834 8188
rect 7770 8128 7834 8132
rect 7850 8188 7914 8192
rect 7850 8132 7854 8188
rect 7854 8132 7910 8188
rect 7910 8132 7914 8188
rect 7850 8128 7914 8132
rect 12049 8188 12113 8192
rect 12049 8132 12053 8188
rect 12053 8132 12109 8188
rect 12109 8132 12113 8188
rect 12049 8128 12113 8132
rect 12129 8188 12193 8192
rect 12129 8132 12133 8188
rect 12133 8132 12189 8188
rect 12189 8132 12193 8188
rect 12129 8128 12193 8132
rect 12209 8188 12273 8192
rect 12209 8132 12213 8188
rect 12213 8132 12269 8188
rect 12269 8132 12273 8188
rect 12209 8128 12273 8132
rect 12289 8188 12353 8192
rect 12289 8132 12293 8188
rect 12293 8132 12349 8188
rect 12349 8132 12353 8188
rect 12289 8128 12353 8132
rect 16488 8188 16552 8192
rect 16488 8132 16492 8188
rect 16492 8132 16548 8188
rect 16548 8132 16552 8188
rect 16488 8128 16552 8132
rect 16568 8188 16632 8192
rect 16568 8132 16572 8188
rect 16572 8132 16628 8188
rect 16628 8132 16632 8188
rect 16568 8128 16632 8132
rect 16648 8188 16712 8192
rect 16648 8132 16652 8188
rect 16652 8132 16708 8188
rect 16708 8132 16712 8188
rect 16648 8128 16712 8132
rect 16728 8188 16792 8192
rect 16728 8132 16732 8188
rect 16732 8132 16788 8188
rect 16788 8132 16792 8188
rect 16728 8128 16792 8132
rect 11284 8060 11348 8124
rect 3831 7644 3895 7648
rect 3831 7588 3835 7644
rect 3835 7588 3891 7644
rect 3891 7588 3895 7644
rect 3831 7584 3895 7588
rect 3911 7644 3975 7648
rect 3911 7588 3915 7644
rect 3915 7588 3971 7644
rect 3971 7588 3975 7644
rect 3911 7584 3975 7588
rect 3991 7644 4055 7648
rect 3991 7588 3995 7644
rect 3995 7588 4051 7644
rect 4051 7588 4055 7644
rect 3991 7584 4055 7588
rect 4071 7644 4135 7648
rect 4071 7588 4075 7644
rect 4075 7588 4131 7644
rect 4131 7588 4135 7644
rect 4071 7584 4135 7588
rect 8270 7644 8334 7648
rect 8270 7588 8274 7644
rect 8274 7588 8330 7644
rect 8330 7588 8334 7644
rect 8270 7584 8334 7588
rect 8350 7644 8414 7648
rect 8350 7588 8354 7644
rect 8354 7588 8410 7644
rect 8410 7588 8414 7644
rect 8350 7584 8414 7588
rect 8430 7644 8494 7648
rect 8430 7588 8434 7644
rect 8434 7588 8490 7644
rect 8490 7588 8494 7644
rect 8430 7584 8494 7588
rect 8510 7644 8574 7648
rect 8510 7588 8514 7644
rect 8514 7588 8570 7644
rect 8570 7588 8574 7644
rect 8510 7584 8574 7588
rect 12709 7644 12773 7648
rect 12709 7588 12713 7644
rect 12713 7588 12769 7644
rect 12769 7588 12773 7644
rect 12709 7584 12773 7588
rect 12789 7644 12853 7648
rect 12789 7588 12793 7644
rect 12793 7588 12849 7644
rect 12849 7588 12853 7644
rect 12789 7584 12853 7588
rect 12869 7644 12933 7648
rect 12869 7588 12873 7644
rect 12873 7588 12929 7644
rect 12929 7588 12933 7644
rect 12869 7584 12933 7588
rect 12949 7644 13013 7648
rect 12949 7588 12953 7644
rect 12953 7588 13009 7644
rect 13009 7588 13013 7644
rect 12949 7584 13013 7588
rect 17148 7644 17212 7648
rect 17148 7588 17152 7644
rect 17152 7588 17208 7644
rect 17208 7588 17212 7644
rect 17148 7584 17212 7588
rect 17228 7644 17292 7648
rect 17228 7588 17232 7644
rect 17232 7588 17288 7644
rect 17288 7588 17292 7644
rect 17228 7584 17292 7588
rect 17308 7644 17372 7648
rect 17308 7588 17312 7644
rect 17312 7588 17368 7644
rect 17368 7588 17372 7644
rect 17308 7584 17372 7588
rect 17388 7644 17452 7648
rect 17388 7588 17392 7644
rect 17392 7588 17448 7644
rect 17448 7588 17452 7644
rect 17388 7584 17452 7588
rect 11652 7516 11716 7580
rect 11836 7516 11900 7580
rect 13492 7516 13556 7580
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 4292 7032 4356 7036
rect 4292 6976 4342 7032
rect 4342 6976 4356 7032
rect 4292 6972 4356 6976
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 13676 6972 13740 7036
rect 14412 6836 14476 6900
rect 1348 6700 1412 6764
rect 11100 6700 11164 6764
rect 11468 6700 11532 6764
rect 3831 6556 3895 6560
rect 3831 6500 3835 6556
rect 3835 6500 3891 6556
rect 3891 6500 3895 6556
rect 3831 6496 3895 6500
rect 3911 6556 3975 6560
rect 3911 6500 3915 6556
rect 3915 6500 3971 6556
rect 3971 6500 3975 6556
rect 3911 6496 3975 6500
rect 3991 6556 4055 6560
rect 3991 6500 3995 6556
rect 3995 6500 4051 6556
rect 4051 6500 4055 6556
rect 3991 6496 4055 6500
rect 4071 6556 4135 6560
rect 4071 6500 4075 6556
rect 4075 6500 4131 6556
rect 4131 6500 4135 6556
rect 4071 6496 4135 6500
rect 8270 6556 8334 6560
rect 8270 6500 8274 6556
rect 8274 6500 8330 6556
rect 8330 6500 8334 6556
rect 8270 6496 8334 6500
rect 8350 6556 8414 6560
rect 8350 6500 8354 6556
rect 8354 6500 8410 6556
rect 8410 6500 8414 6556
rect 8350 6496 8414 6500
rect 8430 6556 8494 6560
rect 8430 6500 8434 6556
rect 8434 6500 8490 6556
rect 8490 6500 8494 6556
rect 8430 6496 8494 6500
rect 8510 6556 8574 6560
rect 8510 6500 8514 6556
rect 8514 6500 8570 6556
rect 8570 6500 8574 6556
rect 8510 6496 8574 6500
rect 12709 6556 12773 6560
rect 12709 6500 12713 6556
rect 12713 6500 12769 6556
rect 12769 6500 12773 6556
rect 12709 6496 12773 6500
rect 12789 6556 12853 6560
rect 12789 6500 12793 6556
rect 12793 6500 12849 6556
rect 12849 6500 12853 6556
rect 12789 6496 12853 6500
rect 12869 6556 12933 6560
rect 12869 6500 12873 6556
rect 12873 6500 12929 6556
rect 12929 6500 12933 6556
rect 12869 6496 12933 6500
rect 12949 6556 13013 6560
rect 12949 6500 12953 6556
rect 12953 6500 13009 6556
rect 13009 6500 13013 6556
rect 12949 6496 13013 6500
rect 17148 6556 17212 6560
rect 17148 6500 17152 6556
rect 17152 6500 17208 6556
rect 17208 6500 17212 6556
rect 17148 6496 17212 6500
rect 17228 6556 17292 6560
rect 17228 6500 17232 6556
rect 17232 6500 17288 6556
rect 17288 6500 17292 6556
rect 17228 6496 17292 6500
rect 17308 6556 17372 6560
rect 17308 6500 17312 6556
rect 17312 6500 17368 6556
rect 17368 6500 17372 6556
rect 17308 6496 17372 6500
rect 17388 6556 17452 6560
rect 17388 6500 17392 6556
rect 17392 6500 17448 6556
rect 17448 6500 17452 6556
rect 17388 6496 17452 6500
rect 9444 6488 9508 6492
rect 9444 6432 9494 6488
rect 9494 6432 9508 6488
rect 9444 6428 9508 6432
rect 11284 6428 11348 6492
rect 10180 6292 10244 6356
rect 17540 6352 17604 6356
rect 17540 6296 17554 6352
rect 17554 6296 17604 6352
rect 6684 6156 6748 6220
rect 17540 6292 17604 6296
rect 12572 6080 12636 6084
rect 12572 6024 12586 6080
rect 12586 6024 12636 6080
rect 12572 6020 12636 6024
rect 13308 6020 13372 6084
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 8892 5884 8956 5948
rect 14596 5884 14660 5948
rect 9812 5748 9876 5812
rect 6684 5612 6748 5676
rect 5396 5476 5460 5540
rect 10548 5536 10612 5540
rect 10548 5480 10598 5536
rect 10598 5480 10612 5536
rect 10548 5476 10612 5480
rect 3831 5468 3895 5472
rect 3831 5412 3835 5468
rect 3835 5412 3891 5468
rect 3891 5412 3895 5468
rect 3831 5408 3895 5412
rect 3911 5468 3975 5472
rect 3911 5412 3915 5468
rect 3915 5412 3971 5468
rect 3971 5412 3975 5468
rect 3911 5408 3975 5412
rect 3991 5468 4055 5472
rect 3991 5412 3995 5468
rect 3995 5412 4051 5468
rect 4051 5412 4055 5468
rect 3991 5408 4055 5412
rect 4071 5468 4135 5472
rect 4071 5412 4075 5468
rect 4075 5412 4131 5468
rect 4131 5412 4135 5468
rect 4071 5408 4135 5412
rect 8270 5468 8334 5472
rect 8270 5412 8274 5468
rect 8274 5412 8330 5468
rect 8330 5412 8334 5468
rect 8270 5408 8334 5412
rect 8350 5468 8414 5472
rect 8350 5412 8354 5468
rect 8354 5412 8410 5468
rect 8410 5412 8414 5468
rect 8350 5408 8414 5412
rect 8430 5468 8494 5472
rect 8430 5412 8434 5468
rect 8434 5412 8490 5468
rect 8490 5412 8494 5468
rect 8430 5408 8494 5412
rect 8510 5468 8574 5472
rect 8510 5412 8514 5468
rect 8514 5412 8570 5468
rect 8570 5412 8574 5468
rect 8510 5408 8574 5412
rect 12709 5468 12773 5472
rect 12709 5412 12713 5468
rect 12713 5412 12769 5468
rect 12769 5412 12773 5468
rect 12709 5408 12773 5412
rect 12789 5468 12853 5472
rect 12789 5412 12793 5468
rect 12793 5412 12849 5468
rect 12849 5412 12853 5468
rect 12789 5408 12853 5412
rect 12869 5468 12933 5472
rect 12869 5412 12873 5468
rect 12873 5412 12929 5468
rect 12929 5412 12933 5468
rect 12869 5408 12933 5412
rect 12949 5468 13013 5472
rect 12949 5412 12953 5468
rect 12953 5412 13009 5468
rect 13009 5412 13013 5468
rect 12949 5408 13013 5412
rect 17148 5468 17212 5472
rect 17148 5412 17152 5468
rect 17152 5412 17208 5468
rect 17208 5412 17212 5468
rect 17148 5408 17212 5412
rect 17228 5468 17292 5472
rect 17228 5412 17232 5468
rect 17232 5412 17288 5468
rect 17288 5412 17292 5468
rect 17228 5408 17292 5412
rect 17308 5468 17372 5472
rect 17308 5412 17312 5468
rect 17312 5412 17368 5468
rect 17368 5412 17372 5468
rect 17308 5408 17372 5412
rect 17388 5468 17452 5472
rect 17388 5412 17392 5468
rect 17392 5412 17448 5468
rect 17448 5412 17452 5468
rect 17388 5408 17452 5412
rect 2636 5204 2700 5268
rect 8708 5204 8772 5268
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5028 4584 5092 4588
rect 5028 4528 5042 4584
rect 5042 4528 5092 4584
rect 5028 4524 5092 4528
rect 6132 4388 6196 4452
rect 3831 4380 3895 4384
rect 3831 4324 3835 4380
rect 3835 4324 3891 4380
rect 3891 4324 3895 4380
rect 3831 4320 3895 4324
rect 3911 4380 3975 4384
rect 3911 4324 3915 4380
rect 3915 4324 3971 4380
rect 3971 4324 3975 4380
rect 3911 4320 3975 4324
rect 3991 4380 4055 4384
rect 3991 4324 3995 4380
rect 3995 4324 4051 4380
rect 4051 4324 4055 4380
rect 3991 4320 4055 4324
rect 4071 4380 4135 4384
rect 4071 4324 4075 4380
rect 4075 4324 4131 4380
rect 4131 4324 4135 4380
rect 4071 4320 4135 4324
rect 8270 4380 8334 4384
rect 8270 4324 8274 4380
rect 8274 4324 8330 4380
rect 8330 4324 8334 4380
rect 8270 4320 8334 4324
rect 8350 4380 8414 4384
rect 8350 4324 8354 4380
rect 8354 4324 8410 4380
rect 8410 4324 8414 4380
rect 8350 4320 8414 4324
rect 8430 4380 8494 4384
rect 8430 4324 8434 4380
rect 8434 4324 8490 4380
rect 8490 4324 8494 4380
rect 8430 4320 8494 4324
rect 8510 4380 8574 4384
rect 8510 4324 8514 4380
rect 8514 4324 8570 4380
rect 8570 4324 8574 4380
rect 8510 4320 8574 4324
rect 3004 4176 3068 4180
rect 3004 4120 3018 4176
rect 3018 4120 3068 4176
rect 3004 4116 3068 4120
rect 9628 4116 9692 4180
rect 12709 4380 12773 4384
rect 12709 4324 12713 4380
rect 12713 4324 12769 4380
rect 12769 4324 12773 4380
rect 12709 4320 12773 4324
rect 12789 4380 12853 4384
rect 12789 4324 12793 4380
rect 12793 4324 12849 4380
rect 12849 4324 12853 4380
rect 12789 4320 12853 4324
rect 12869 4380 12933 4384
rect 12869 4324 12873 4380
rect 12873 4324 12929 4380
rect 12929 4324 12933 4380
rect 12869 4320 12933 4324
rect 12949 4380 13013 4384
rect 12949 4324 12953 4380
rect 12953 4324 13009 4380
rect 13009 4324 13013 4380
rect 12949 4320 13013 4324
rect 17148 4380 17212 4384
rect 17148 4324 17152 4380
rect 17152 4324 17208 4380
rect 17208 4324 17212 4380
rect 17148 4320 17212 4324
rect 17228 4380 17292 4384
rect 17228 4324 17232 4380
rect 17232 4324 17288 4380
rect 17288 4324 17292 4380
rect 17228 4320 17292 4324
rect 17308 4380 17372 4384
rect 17308 4324 17312 4380
rect 17312 4324 17368 4380
rect 17368 4324 17372 4380
rect 17308 4320 17372 4324
rect 17388 4380 17452 4384
rect 17388 4324 17392 4380
rect 17392 4324 17448 4380
rect 17448 4324 17452 4380
rect 17388 4320 17452 4324
rect 1164 3980 1228 4044
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 796 3708 860 3772
rect 6500 3768 6564 3772
rect 6500 3712 6514 3768
rect 6514 3712 6564 3768
rect 6500 3708 6564 3712
rect 15516 3768 15580 3772
rect 15516 3712 15530 3768
rect 15530 3712 15580 3768
rect 15516 3708 15580 3712
rect 15148 3436 15212 3500
rect 3831 3292 3895 3296
rect 3831 3236 3835 3292
rect 3835 3236 3891 3292
rect 3891 3236 3895 3292
rect 3831 3232 3895 3236
rect 3911 3292 3975 3296
rect 3911 3236 3915 3292
rect 3915 3236 3971 3292
rect 3971 3236 3975 3292
rect 3911 3232 3975 3236
rect 3991 3292 4055 3296
rect 3991 3236 3995 3292
rect 3995 3236 4051 3292
rect 4051 3236 4055 3292
rect 3991 3232 4055 3236
rect 4071 3292 4135 3296
rect 4071 3236 4075 3292
rect 4075 3236 4131 3292
rect 4131 3236 4135 3292
rect 4071 3232 4135 3236
rect 8270 3292 8334 3296
rect 8270 3236 8274 3292
rect 8274 3236 8330 3292
rect 8330 3236 8334 3292
rect 8270 3232 8334 3236
rect 8350 3292 8414 3296
rect 8350 3236 8354 3292
rect 8354 3236 8410 3292
rect 8410 3236 8414 3292
rect 8350 3232 8414 3236
rect 8430 3292 8494 3296
rect 8430 3236 8434 3292
rect 8434 3236 8490 3292
rect 8490 3236 8494 3292
rect 8430 3232 8494 3236
rect 8510 3292 8574 3296
rect 8510 3236 8514 3292
rect 8514 3236 8570 3292
rect 8570 3236 8574 3292
rect 8510 3232 8574 3236
rect 12709 3292 12773 3296
rect 12709 3236 12713 3292
rect 12713 3236 12769 3292
rect 12769 3236 12773 3292
rect 12709 3232 12773 3236
rect 12789 3292 12853 3296
rect 12789 3236 12793 3292
rect 12793 3236 12849 3292
rect 12849 3236 12853 3292
rect 12789 3232 12853 3236
rect 12869 3292 12933 3296
rect 12869 3236 12873 3292
rect 12873 3236 12929 3292
rect 12929 3236 12933 3292
rect 12869 3232 12933 3236
rect 12949 3292 13013 3296
rect 12949 3236 12953 3292
rect 12953 3236 13009 3292
rect 13009 3236 13013 3292
rect 12949 3232 13013 3236
rect 17148 3292 17212 3296
rect 17148 3236 17152 3292
rect 17152 3236 17208 3292
rect 17208 3236 17212 3292
rect 17148 3232 17212 3236
rect 17228 3292 17292 3296
rect 17228 3236 17232 3292
rect 17232 3236 17288 3292
rect 17288 3236 17292 3292
rect 17228 3232 17292 3236
rect 17308 3292 17372 3296
rect 17308 3236 17312 3292
rect 17312 3236 17368 3292
rect 17368 3236 17372 3292
rect 17308 3232 17372 3236
rect 17388 3292 17452 3296
rect 17388 3236 17392 3292
rect 17392 3236 17448 3292
rect 17448 3236 17452 3292
rect 17388 3232 17452 3236
rect 17908 3164 17972 3228
rect 980 3028 1044 3092
rect 14964 2892 15028 2956
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 3831 2204 3895 2208
rect 3831 2148 3835 2204
rect 3835 2148 3891 2204
rect 3891 2148 3895 2204
rect 3831 2144 3895 2148
rect 3911 2204 3975 2208
rect 3911 2148 3915 2204
rect 3915 2148 3971 2204
rect 3971 2148 3975 2204
rect 3911 2144 3975 2148
rect 3991 2204 4055 2208
rect 3991 2148 3995 2204
rect 3995 2148 4051 2204
rect 4051 2148 4055 2204
rect 3991 2144 4055 2148
rect 4071 2204 4135 2208
rect 4071 2148 4075 2204
rect 4075 2148 4131 2204
rect 4131 2148 4135 2204
rect 4071 2144 4135 2148
rect 8270 2204 8334 2208
rect 8270 2148 8274 2204
rect 8274 2148 8330 2204
rect 8330 2148 8334 2204
rect 8270 2144 8334 2148
rect 8350 2204 8414 2208
rect 8350 2148 8354 2204
rect 8354 2148 8410 2204
rect 8410 2148 8414 2204
rect 8350 2144 8414 2148
rect 8430 2204 8494 2208
rect 8430 2148 8434 2204
rect 8434 2148 8490 2204
rect 8490 2148 8494 2204
rect 8430 2144 8494 2148
rect 8510 2204 8574 2208
rect 8510 2148 8514 2204
rect 8514 2148 8570 2204
rect 8570 2148 8574 2204
rect 8510 2144 8574 2148
rect 12709 2204 12773 2208
rect 12709 2148 12713 2204
rect 12713 2148 12769 2204
rect 12769 2148 12773 2204
rect 12709 2144 12773 2148
rect 12789 2204 12853 2208
rect 12789 2148 12793 2204
rect 12793 2148 12849 2204
rect 12849 2148 12853 2204
rect 12789 2144 12853 2148
rect 12869 2204 12933 2208
rect 12869 2148 12873 2204
rect 12873 2148 12929 2204
rect 12929 2148 12933 2204
rect 12869 2144 12933 2148
rect 12949 2204 13013 2208
rect 12949 2148 12953 2204
rect 12953 2148 13009 2204
rect 13009 2148 13013 2204
rect 12949 2144 13013 2148
rect 17148 2204 17212 2208
rect 17148 2148 17152 2204
rect 17152 2148 17208 2204
rect 17208 2148 17212 2204
rect 17148 2144 17212 2148
rect 17228 2204 17292 2208
rect 17228 2148 17232 2204
rect 17232 2148 17288 2204
rect 17288 2148 17292 2204
rect 17228 2144 17292 2148
rect 17308 2204 17372 2208
rect 17308 2148 17312 2204
rect 17312 2148 17368 2204
rect 17368 2148 17372 2204
rect 17308 2144 17372 2148
rect 17388 2204 17452 2208
rect 17388 2148 17392 2204
rect 17392 2148 17448 2204
rect 17448 2148 17452 2204
rect 17388 2144 17452 2148
<< metal4 >>
rect 9259 19820 9325 19821
rect 9259 19756 9260 19820
rect 9324 19756 9325 19820
rect 9259 19755 9325 19756
rect -1076 19546 -756 19588
rect -1076 19310 -1034 19546
rect -798 19310 -756 19546
rect -1076 16282 -756 19310
rect -1076 16046 -1034 16282
rect -798 16046 -756 16282
rect -1076 12474 -756 16046
rect -1076 12238 -1034 12474
rect -798 12238 -756 12474
rect -1076 8666 -756 12238
rect -1076 8430 -1034 8666
rect -798 8430 -756 8666
rect -1076 4858 -756 8430
rect -1076 4622 -1034 4858
rect -798 4622 -756 4858
rect -1076 274 -756 4622
rect -416 18886 -96 18928
rect -416 18650 -374 18886
rect -138 18650 -96 18886
rect -416 15622 -96 18650
rect 3163 18886 3483 19588
rect 3163 18650 3205 18886
rect 3441 18650 3483 18886
rect 1347 18052 1413 18053
rect 1347 17988 1348 18052
rect 1412 17988 1413 18052
rect 1347 17987 1413 17988
rect 1163 17644 1229 17645
rect 1163 17580 1164 17644
rect 1228 17580 1229 17644
rect 1163 17579 1229 17580
rect -416 15386 -374 15622
rect -138 15386 -96 15622
rect -416 11814 -96 15386
rect 795 14108 861 14109
rect 795 14044 796 14108
rect 860 14044 861 14108
rect 795 14043 861 14044
rect -416 11578 -374 11814
rect -138 11578 -96 11814
rect -416 8006 -96 11578
rect -416 7770 -374 8006
rect -138 7770 -96 8006
rect -416 4198 -96 7770
rect -416 3962 -374 4198
rect -138 3962 -96 4198
rect -416 934 -96 3962
rect 798 3773 858 14043
rect 979 13836 1045 13837
rect 979 13772 980 13836
rect 1044 13772 1045 13836
rect 979 13771 1045 13772
rect 795 3772 861 3773
rect 795 3708 796 3772
rect 860 3708 861 3772
rect 795 3707 861 3708
rect 982 3093 1042 13771
rect 1166 4045 1226 17579
rect 1350 6765 1410 17987
rect 3163 16896 3483 18650
rect 3163 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3483 16896
rect 3003 16692 3069 16693
rect 3003 16628 3004 16692
rect 3068 16628 3069 16692
rect 3003 16627 3069 16628
rect 2635 16556 2701 16557
rect 2635 16492 2636 16556
rect 2700 16492 2701 16556
rect 2635 16491 2701 16492
rect 1347 6764 1413 6765
rect 1347 6700 1348 6764
rect 1412 6700 1413 6764
rect 1347 6699 1413 6700
rect 2638 5269 2698 16491
rect 2635 5268 2701 5269
rect 2635 5204 2636 5268
rect 2700 5204 2701 5268
rect 2635 5203 2701 5204
rect 3006 4181 3066 16627
rect 3163 15808 3483 16832
rect 3823 19546 4143 19588
rect 3823 19310 3865 19546
rect 4101 19310 4143 19546
rect 3823 17440 4143 19310
rect 3823 17376 3831 17440
rect 3895 17376 3911 17440
rect 3975 17376 3991 17440
rect 4055 17376 4071 17440
rect 4135 17376 4143 17440
rect 3823 16352 4143 17376
rect 3823 16288 3831 16352
rect 3895 16288 3911 16352
rect 3975 16288 3991 16352
rect 4055 16288 4071 16352
rect 4135 16288 4143 16352
rect 3823 16282 4143 16288
rect 7602 18886 7922 19588
rect 7602 18650 7644 18886
rect 7880 18650 7922 18886
rect 7602 16896 7922 18650
rect 7602 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7922 16896
rect 3555 16148 3621 16149
rect 3555 16084 3556 16148
rect 3620 16084 3621 16148
rect 3555 16083 3621 16084
rect 3163 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3483 15808
rect 3163 15622 3483 15744
rect 3163 15386 3205 15622
rect 3441 15386 3483 15622
rect 3163 14720 3483 15386
rect 3163 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3483 14720
rect 3163 13632 3483 14656
rect 3163 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3483 13632
rect 3163 12544 3483 13568
rect 3558 12749 3618 16083
rect 3823 16046 3865 16282
rect 4101 16046 4143 16282
rect 4475 16284 4541 16285
rect 4475 16220 4476 16284
rect 4540 16220 4541 16284
rect 4475 16219 4541 16220
rect 3823 15264 4143 16046
rect 3823 15200 3831 15264
rect 3895 15200 3911 15264
rect 3975 15200 3991 15264
rect 4055 15200 4071 15264
rect 4135 15200 4143 15264
rect 3823 14176 4143 15200
rect 3823 14112 3831 14176
rect 3895 14112 3911 14176
rect 3975 14112 3991 14176
rect 4055 14112 4071 14176
rect 4135 14112 4143 14176
rect 3823 13088 4143 14112
rect 4291 14108 4357 14109
rect 4291 14044 4292 14108
rect 4356 14044 4357 14108
rect 4291 14043 4357 14044
rect 3823 13024 3831 13088
rect 3895 13024 3911 13088
rect 3975 13024 3991 13088
rect 4055 13024 4071 13088
rect 4135 13024 4143 13088
rect 3555 12748 3621 12749
rect 3555 12684 3556 12748
rect 3620 12684 3621 12748
rect 3555 12683 3621 12684
rect 3163 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3483 12544
rect 3163 11814 3483 12480
rect 3163 11578 3205 11814
rect 3441 11578 3483 11814
rect 3163 11456 3483 11578
rect 3163 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3483 11456
rect 3163 10368 3483 11392
rect 3163 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3483 10368
rect 3163 9280 3483 10304
rect 3558 9621 3618 12683
rect 3823 12474 4143 13024
rect 3823 12238 3865 12474
rect 4101 12238 4143 12474
rect 4294 12341 4354 14043
rect 4291 12340 4357 12341
rect 4291 12276 4292 12340
rect 4356 12276 4357 12340
rect 4291 12275 4357 12276
rect 3823 12000 4143 12238
rect 3823 11936 3831 12000
rect 3895 11936 3911 12000
rect 3975 11936 3991 12000
rect 4055 11936 4071 12000
rect 4135 11936 4143 12000
rect 3823 10912 4143 11936
rect 3823 10848 3831 10912
rect 3895 10848 3911 10912
rect 3975 10848 3991 10912
rect 4055 10848 4071 10912
rect 4135 10848 4143 10912
rect 3823 9824 4143 10848
rect 4291 10572 4357 10573
rect 4291 10508 4292 10572
rect 4356 10508 4357 10572
rect 4291 10507 4357 10508
rect 3823 9760 3831 9824
rect 3895 9760 3911 9824
rect 3975 9760 3991 9824
rect 4055 9760 4071 9824
rect 4135 9760 4143 9824
rect 3555 9620 3621 9621
rect 3555 9556 3556 9620
rect 3620 9556 3621 9620
rect 3555 9555 3621 9556
rect 3163 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3483 9280
rect 3163 8192 3483 9216
rect 3163 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3483 8192
rect 3163 8006 3483 8128
rect 3163 7770 3205 8006
rect 3441 7770 3483 8006
rect 3163 7104 3483 7770
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 4198 3483 4864
rect 3003 4180 3069 4181
rect 3003 4116 3004 4180
rect 3068 4116 3069 4180
rect 3003 4115 3069 4116
rect 1163 4044 1229 4045
rect 1163 3980 1164 4044
rect 1228 3980 1229 4044
rect 1163 3979 1229 3980
rect 3163 3962 3205 4198
rect 3441 3962 3483 4198
rect 3163 3840 3483 3962
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 979 3092 1045 3093
rect 979 3028 980 3092
rect 1044 3028 1045 3092
rect 979 3027 1045 3028
rect -416 698 -374 934
rect -138 698 -96 934
rect -416 656 -96 698
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 934 3483 2688
rect 3163 698 3205 934
rect 3441 698 3483 934
rect -1076 38 -1034 274
rect -798 38 -756 274
rect -1076 -4 -756 38
rect 3163 -4 3483 698
rect 3823 8736 4143 9760
rect 3823 8672 3831 8736
rect 3895 8672 3911 8736
rect 3975 8672 3991 8736
rect 4055 8672 4071 8736
rect 4135 8672 4143 8736
rect 3823 8666 4143 8672
rect 3823 8430 3865 8666
rect 4101 8430 4143 8666
rect 3823 7648 4143 8430
rect 3823 7584 3831 7648
rect 3895 7584 3911 7648
rect 3975 7584 3991 7648
rect 4055 7584 4071 7648
rect 4135 7584 4143 7648
rect 3823 6560 4143 7584
rect 4294 7037 4354 10507
rect 4478 10437 4538 16219
rect 6867 15876 6933 15877
rect 6867 15812 6868 15876
rect 6932 15812 6933 15876
rect 6867 15811 6933 15812
rect 4843 14108 4909 14109
rect 4843 14044 4844 14108
rect 4908 14044 4909 14108
rect 4843 14043 4909 14044
rect 4846 11253 4906 14043
rect 6499 13564 6565 13565
rect 6499 13500 6500 13564
rect 6564 13500 6565 13564
rect 6499 13499 6565 13500
rect 6131 12612 6197 12613
rect 6131 12548 6132 12612
rect 6196 12548 6197 12612
rect 6131 12547 6197 12548
rect 5027 12476 5093 12477
rect 5027 12412 5028 12476
rect 5092 12412 5093 12476
rect 5027 12411 5093 12412
rect 4843 11252 4909 11253
rect 4843 11188 4844 11252
rect 4908 11188 4909 11252
rect 4843 11187 4909 11188
rect 4475 10436 4541 10437
rect 4475 10372 4476 10436
rect 4540 10372 4541 10436
rect 4475 10371 4541 10372
rect 4291 7036 4357 7037
rect 4291 6972 4292 7036
rect 4356 6972 4357 7036
rect 4291 6971 4357 6972
rect 3823 6496 3831 6560
rect 3895 6496 3911 6560
rect 3975 6496 3991 6560
rect 4055 6496 4071 6560
rect 4135 6496 4143 6560
rect 3823 5472 4143 6496
rect 3823 5408 3831 5472
rect 3895 5408 3911 5472
rect 3975 5408 3991 5472
rect 4055 5408 4071 5472
rect 4135 5408 4143 5472
rect 3823 4858 4143 5408
rect 3823 4622 3865 4858
rect 4101 4622 4143 4858
rect 3823 4384 4143 4622
rect 5030 4589 5090 12411
rect 5395 10708 5461 10709
rect 5395 10644 5396 10708
rect 5460 10644 5461 10708
rect 5395 10643 5461 10644
rect 5398 8805 5458 10643
rect 5395 8804 5461 8805
rect 5395 8740 5396 8804
rect 5460 8740 5461 8804
rect 5395 8739 5461 8740
rect 5398 5541 5458 8739
rect 5395 5540 5461 5541
rect 5395 5476 5396 5540
rect 5460 5476 5461 5540
rect 5395 5475 5461 5476
rect 5027 4588 5093 4589
rect 5027 4524 5028 4588
rect 5092 4524 5093 4588
rect 5027 4523 5093 4524
rect 6134 4453 6194 12547
rect 6315 9484 6381 9485
rect 6315 9420 6316 9484
rect 6380 9420 6381 9484
rect 6315 9419 6381 9420
rect 6318 8669 6378 9419
rect 6502 9077 6562 13499
rect 6683 12068 6749 12069
rect 6683 12004 6684 12068
rect 6748 12004 6749 12068
rect 6683 12003 6749 12004
rect 6499 9076 6565 9077
rect 6499 9012 6500 9076
rect 6564 9012 6565 9076
rect 6499 9011 6565 9012
rect 6315 8668 6381 8669
rect 6315 8604 6316 8668
rect 6380 8604 6381 8668
rect 6315 8603 6381 8604
rect 6131 4452 6197 4453
rect 6131 4388 6132 4452
rect 6196 4388 6197 4452
rect 6131 4387 6197 4388
rect 3823 4320 3831 4384
rect 3895 4320 3911 4384
rect 3975 4320 3991 4384
rect 4055 4320 4071 4384
rect 4135 4320 4143 4384
rect 3823 3296 4143 4320
rect 6502 3773 6562 9011
rect 6686 6221 6746 12003
rect 6870 10437 6930 15811
rect 7602 15808 7922 16832
rect 7602 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7922 15808
rect 7602 15622 7922 15744
rect 7602 15386 7644 15622
rect 7880 15386 7922 15622
rect 7051 15196 7117 15197
rect 7051 15132 7052 15196
rect 7116 15132 7117 15196
rect 7051 15131 7117 15132
rect 6867 10436 6933 10437
rect 6867 10372 6868 10436
rect 6932 10372 6933 10436
rect 6867 10371 6933 10372
rect 7054 10301 7114 15131
rect 7602 14720 7922 15386
rect 7602 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7922 14720
rect 7602 13632 7922 14656
rect 7602 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7922 13632
rect 7235 13156 7301 13157
rect 7235 13092 7236 13156
rect 7300 13092 7301 13156
rect 7235 13091 7301 13092
rect 7051 10300 7117 10301
rect 7051 10236 7052 10300
rect 7116 10236 7117 10300
rect 7051 10235 7117 10236
rect 7238 8941 7298 13091
rect 7602 12544 7922 13568
rect 7602 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7922 12544
rect 7419 11932 7485 11933
rect 7419 11868 7420 11932
rect 7484 11868 7485 11932
rect 7419 11867 7485 11868
rect 7235 8940 7301 8941
rect 7235 8876 7236 8940
rect 7300 8876 7301 8940
rect 7235 8875 7301 8876
rect 7422 8669 7482 11867
rect 7602 11814 7922 12480
rect 7602 11578 7644 11814
rect 7880 11578 7922 11814
rect 7602 11456 7922 11578
rect 7602 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7922 11456
rect 7602 10368 7922 11392
rect 7602 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7922 10368
rect 7602 9280 7922 10304
rect 7602 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7922 9280
rect 7419 8668 7485 8669
rect 7419 8604 7420 8668
rect 7484 8604 7485 8668
rect 7419 8603 7485 8604
rect 7602 8192 7922 9216
rect 7602 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7922 8192
rect 7602 8006 7922 8128
rect 7602 7770 7644 8006
rect 7880 7770 7922 8006
rect 7602 7104 7922 7770
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 6683 6220 6749 6221
rect 6683 6156 6684 6220
rect 6748 6156 6749 6220
rect 6683 6155 6749 6156
rect 6686 5677 6746 6155
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 6683 5676 6749 5677
rect 6683 5612 6684 5676
rect 6748 5612 6749 5676
rect 6683 5611 6749 5612
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 4198 7922 4864
rect 7602 3962 7644 4198
rect 7880 3962 7922 4198
rect 7602 3840 7922 3962
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 6499 3772 6565 3773
rect 6499 3708 6500 3772
rect 6564 3708 6565 3772
rect 6499 3707 6565 3708
rect 3823 3232 3831 3296
rect 3895 3232 3911 3296
rect 3975 3232 3991 3296
rect 4055 3232 4071 3296
rect 4135 3232 4143 3296
rect 3823 2208 4143 3232
rect 3823 2144 3831 2208
rect 3895 2144 3911 2208
rect 3975 2144 3991 2208
rect 4055 2144 4071 2208
rect 4135 2144 4143 2208
rect 3823 274 4143 2144
rect 3823 38 3865 274
rect 4101 38 4143 274
rect 3823 -4 4143 38
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 934 7922 2688
rect 7602 698 7644 934
rect 7880 698 7922 934
rect 7602 -4 7922 698
rect 8262 19546 8582 19588
rect 8262 19310 8304 19546
rect 8540 19310 8582 19546
rect 8262 17440 8582 19310
rect 8262 17376 8270 17440
rect 8334 17376 8350 17440
rect 8414 17376 8430 17440
rect 8494 17376 8510 17440
rect 8574 17376 8582 17440
rect 8262 16352 8582 17376
rect 9075 16964 9141 16965
rect 9075 16900 9076 16964
rect 9140 16900 9141 16964
rect 9075 16899 9141 16900
rect 8262 16288 8270 16352
rect 8334 16288 8350 16352
rect 8414 16288 8430 16352
rect 8494 16288 8510 16352
rect 8574 16288 8582 16352
rect 8262 16282 8582 16288
rect 8262 16046 8304 16282
rect 8540 16046 8582 16282
rect 8262 15264 8582 16046
rect 8262 15200 8270 15264
rect 8334 15200 8350 15264
rect 8414 15200 8430 15264
rect 8494 15200 8510 15264
rect 8574 15200 8582 15264
rect 8262 14176 8582 15200
rect 8707 14788 8773 14789
rect 8707 14724 8708 14788
rect 8772 14724 8773 14788
rect 8707 14723 8773 14724
rect 8262 14112 8270 14176
rect 8334 14112 8350 14176
rect 8414 14112 8430 14176
rect 8494 14112 8510 14176
rect 8574 14112 8582 14176
rect 8262 13088 8582 14112
rect 8262 13024 8270 13088
rect 8334 13024 8350 13088
rect 8414 13024 8430 13088
rect 8494 13024 8510 13088
rect 8574 13024 8582 13088
rect 8262 12474 8582 13024
rect 8262 12238 8304 12474
rect 8540 12238 8582 12474
rect 8710 12341 8770 14723
rect 8707 12340 8773 12341
rect 8707 12276 8708 12340
rect 8772 12276 8773 12340
rect 8707 12275 8773 12276
rect 8262 12000 8582 12238
rect 8262 11936 8270 12000
rect 8334 11936 8350 12000
rect 8414 11936 8430 12000
rect 8494 11936 8510 12000
rect 8574 11936 8582 12000
rect 8262 10912 8582 11936
rect 8891 11660 8957 11661
rect 8891 11596 8892 11660
rect 8956 11596 8957 11660
rect 8891 11595 8957 11596
rect 8707 10980 8773 10981
rect 8707 10916 8708 10980
rect 8772 10916 8773 10980
rect 8707 10915 8773 10916
rect 8262 10848 8270 10912
rect 8334 10848 8350 10912
rect 8414 10848 8430 10912
rect 8494 10848 8510 10912
rect 8574 10848 8582 10912
rect 8262 9824 8582 10848
rect 8710 10437 8770 10915
rect 8707 10436 8773 10437
rect 8707 10372 8708 10436
rect 8772 10372 8773 10436
rect 8707 10371 8773 10372
rect 8262 9760 8270 9824
rect 8334 9760 8350 9824
rect 8414 9760 8430 9824
rect 8494 9760 8510 9824
rect 8574 9760 8582 9824
rect 8262 8736 8582 9760
rect 8262 8672 8270 8736
rect 8334 8672 8350 8736
rect 8414 8672 8430 8736
rect 8494 8672 8510 8736
rect 8574 8672 8582 8736
rect 8262 8666 8582 8672
rect 8262 8430 8304 8666
rect 8540 8430 8582 8666
rect 8262 7648 8582 8430
rect 8262 7584 8270 7648
rect 8334 7584 8350 7648
rect 8414 7584 8430 7648
rect 8494 7584 8510 7648
rect 8574 7584 8582 7648
rect 8262 6560 8582 7584
rect 8262 6496 8270 6560
rect 8334 6496 8350 6560
rect 8414 6496 8430 6560
rect 8494 6496 8510 6560
rect 8574 6496 8582 6560
rect 8262 5472 8582 6496
rect 8262 5408 8270 5472
rect 8334 5408 8350 5472
rect 8414 5408 8430 5472
rect 8494 5408 8510 5472
rect 8574 5408 8582 5472
rect 8262 4858 8582 5408
rect 8710 5269 8770 10371
rect 8894 5949 8954 11595
rect 9078 10709 9138 16899
rect 9075 10708 9141 10709
rect 9075 10644 9076 10708
rect 9140 10644 9141 10708
rect 9075 10643 9141 10644
rect 9262 10301 9322 19755
rect 12041 18886 12361 19588
rect 12041 18650 12083 18886
rect 12319 18650 12361 18886
rect 12041 16896 12361 18650
rect 12041 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12361 16896
rect 9627 16828 9693 16829
rect 9627 16764 9628 16828
rect 9692 16764 9693 16828
rect 9627 16763 9693 16764
rect 9443 13292 9509 13293
rect 9443 13228 9444 13292
rect 9508 13228 9509 13292
rect 9443 13227 9509 13228
rect 9446 10437 9506 13227
rect 9443 10436 9509 10437
rect 9443 10372 9444 10436
rect 9508 10372 9509 10436
rect 9443 10371 9509 10372
rect 9259 10300 9325 10301
rect 9259 10236 9260 10300
rect 9324 10236 9325 10300
rect 9259 10235 9325 10236
rect 9446 6493 9506 10371
rect 9443 6492 9509 6493
rect 9443 6428 9444 6492
rect 9508 6428 9509 6492
rect 9443 6427 9509 6428
rect 8891 5948 8957 5949
rect 8891 5884 8892 5948
rect 8956 5884 8957 5948
rect 8891 5883 8957 5884
rect 8707 5268 8773 5269
rect 8707 5204 8708 5268
rect 8772 5204 8773 5268
rect 8707 5203 8773 5204
rect 8262 4622 8304 4858
rect 8540 4622 8582 4858
rect 8262 4384 8582 4622
rect 8262 4320 8270 4384
rect 8334 4320 8350 4384
rect 8414 4320 8430 4384
rect 8494 4320 8510 4384
rect 8574 4320 8582 4384
rect 8262 3296 8582 4320
rect 9630 4181 9690 16763
rect 9995 16284 10061 16285
rect 9995 16220 9996 16284
rect 10060 16220 10061 16284
rect 9995 16219 10061 16220
rect 9811 13156 9877 13157
rect 9811 13092 9812 13156
rect 9876 13092 9877 13156
rect 9811 13091 9877 13092
rect 9814 12613 9874 13091
rect 9811 12612 9877 12613
rect 9811 12548 9812 12612
rect 9876 12548 9877 12612
rect 9811 12547 9877 12548
rect 9811 12340 9877 12341
rect 9811 12276 9812 12340
rect 9876 12276 9877 12340
rect 9811 12275 9877 12276
rect 9814 11933 9874 12275
rect 9811 11932 9877 11933
rect 9811 11868 9812 11932
rect 9876 11868 9877 11932
rect 9811 11867 9877 11868
rect 9814 10301 9874 11867
rect 9811 10300 9877 10301
rect 9811 10236 9812 10300
rect 9876 10236 9877 10300
rect 9811 10235 9877 10236
rect 9811 9756 9877 9757
rect 9811 9692 9812 9756
rect 9876 9692 9877 9756
rect 9811 9691 9877 9692
rect 9814 5813 9874 9691
rect 9998 8261 10058 16219
rect 12041 15808 12361 16832
rect 12041 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12361 15808
rect 12041 15622 12361 15744
rect 12041 15386 12083 15622
rect 12319 15386 12361 15622
rect 12041 14720 12361 15386
rect 12041 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12361 14720
rect 11467 14652 11533 14653
rect 11467 14588 11468 14652
rect 11532 14588 11533 14652
rect 11467 14587 11533 14588
rect 11099 14516 11165 14517
rect 11099 14452 11100 14516
rect 11164 14452 11165 14516
rect 11099 14451 11165 14452
rect 10731 14244 10797 14245
rect 10731 14180 10732 14244
rect 10796 14180 10797 14244
rect 10731 14179 10797 14180
rect 10363 13972 10429 13973
rect 10363 13908 10364 13972
rect 10428 13908 10429 13972
rect 10363 13907 10429 13908
rect 10179 11932 10245 11933
rect 10179 11868 10180 11932
rect 10244 11868 10245 11932
rect 10179 11867 10245 11868
rect 9995 8260 10061 8261
rect 9995 8196 9996 8260
rect 10060 8196 10061 8260
rect 9995 8195 10061 8196
rect 10182 6357 10242 11867
rect 10366 10709 10426 13907
rect 10734 11525 10794 14179
rect 10731 11524 10797 11525
rect 10731 11460 10732 11524
rect 10796 11460 10797 11524
rect 10731 11459 10797 11460
rect 10547 11388 10613 11389
rect 10547 11324 10548 11388
rect 10612 11324 10613 11388
rect 10547 11323 10613 11324
rect 10363 10708 10429 10709
rect 10363 10644 10364 10708
rect 10428 10644 10429 10708
rect 10363 10643 10429 10644
rect 10179 6356 10245 6357
rect 10179 6292 10180 6356
rect 10244 6292 10245 6356
rect 10179 6291 10245 6292
rect 9811 5812 9877 5813
rect 9811 5748 9812 5812
rect 9876 5748 9877 5812
rect 9811 5747 9877 5748
rect 10550 5541 10610 11323
rect 11102 10709 11162 14451
rect 11099 10708 11165 10709
rect 11099 10644 11100 10708
rect 11164 10644 11165 10708
rect 11099 10643 11165 10644
rect 11099 8396 11165 8397
rect 11099 8332 11100 8396
rect 11164 8332 11165 8396
rect 11099 8331 11165 8332
rect 11102 6765 11162 8331
rect 11283 8124 11349 8125
rect 11283 8060 11284 8124
rect 11348 8060 11349 8124
rect 11283 8059 11349 8060
rect 11099 6764 11165 6765
rect 11099 6700 11100 6764
rect 11164 6700 11165 6764
rect 11099 6699 11165 6700
rect 11286 6493 11346 8059
rect 11470 6765 11530 14587
rect 11835 13700 11901 13701
rect 11835 13636 11836 13700
rect 11900 13636 11901 13700
rect 11835 13635 11901 13636
rect 11651 12204 11717 12205
rect 11651 12140 11652 12204
rect 11716 12140 11717 12204
rect 11651 12139 11717 12140
rect 11654 9621 11714 12139
rect 11838 10709 11898 13635
rect 12041 13632 12361 14656
rect 12041 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12361 13632
rect 12041 12544 12361 13568
rect 12041 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12361 12544
rect 12041 11814 12361 12480
rect 12041 11578 12083 11814
rect 12319 11578 12361 11814
rect 12041 11456 12361 11578
rect 12041 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12361 11456
rect 11835 10708 11901 10709
rect 11835 10644 11836 10708
rect 11900 10644 11901 10708
rect 11835 10643 11901 10644
rect 12041 10368 12361 11392
rect 12041 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12361 10368
rect 11835 10164 11901 10165
rect 11835 10100 11836 10164
rect 11900 10100 11901 10164
rect 11835 10099 11901 10100
rect 11651 9620 11717 9621
rect 11651 9556 11652 9620
rect 11716 9556 11717 9620
rect 11651 9555 11717 9556
rect 11651 9212 11717 9213
rect 11651 9148 11652 9212
rect 11716 9148 11717 9212
rect 11651 9147 11717 9148
rect 11654 7581 11714 9147
rect 11838 7581 11898 10099
rect 12041 9280 12361 10304
rect 12701 19546 13021 19588
rect 12701 19310 12743 19546
rect 12979 19310 13021 19546
rect 12701 17440 13021 19310
rect 12701 17376 12709 17440
rect 12773 17376 12789 17440
rect 12853 17376 12869 17440
rect 12933 17376 12949 17440
rect 13013 17376 13021 17440
rect 12701 16352 13021 17376
rect 12701 16288 12709 16352
rect 12773 16288 12789 16352
rect 12853 16288 12869 16352
rect 12933 16288 12949 16352
rect 13013 16288 13021 16352
rect 12701 16282 13021 16288
rect 12701 16046 12743 16282
rect 12979 16046 13021 16282
rect 12701 15264 13021 16046
rect 16480 18886 16800 19588
rect 16480 18650 16522 18886
rect 16758 18650 16800 18886
rect 16480 16896 16800 18650
rect 17140 19546 17460 19588
rect 17140 19310 17182 19546
rect 17418 19310 17460 19546
rect 16987 18188 17053 18189
rect 16987 18124 16988 18188
rect 17052 18124 17053 18188
rect 16987 18123 17053 18124
rect 16480 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16800 16896
rect 14779 16012 14845 16013
rect 14779 15948 14780 16012
rect 14844 15948 14845 16012
rect 14779 15947 14845 15948
rect 14595 15332 14661 15333
rect 14595 15268 14596 15332
rect 14660 15268 14661 15332
rect 14595 15267 14661 15268
rect 12701 15200 12709 15264
rect 12773 15200 12789 15264
rect 12853 15200 12869 15264
rect 12933 15200 12949 15264
rect 13013 15200 13021 15264
rect 12701 14176 13021 15200
rect 12701 14112 12709 14176
rect 12773 14112 12789 14176
rect 12853 14112 12869 14176
rect 12933 14112 12949 14176
rect 13013 14112 13021 14176
rect 12701 13088 13021 14112
rect 13307 13836 13373 13837
rect 13307 13772 13308 13836
rect 13372 13772 13373 13836
rect 13307 13771 13373 13772
rect 12701 13024 12709 13088
rect 12773 13024 12789 13088
rect 12853 13024 12869 13088
rect 12933 13024 12949 13088
rect 13013 13024 13021 13088
rect 12701 12474 13021 13024
rect 12701 12238 12743 12474
rect 12979 12238 13021 12474
rect 12701 12000 13021 12238
rect 12701 11936 12709 12000
rect 12773 11936 12789 12000
rect 12853 11936 12869 12000
rect 12933 11936 12949 12000
rect 13013 11936 13021 12000
rect 12701 10912 13021 11936
rect 12701 10848 12709 10912
rect 12773 10848 12789 10912
rect 12853 10848 12869 10912
rect 12933 10848 12949 10912
rect 13013 10848 13021 10912
rect 12701 9824 13021 10848
rect 12701 9760 12709 9824
rect 12773 9760 12789 9824
rect 12853 9760 12869 9824
rect 12933 9760 12949 9824
rect 13013 9760 13021 9824
rect 12571 9348 12637 9349
rect 12571 9284 12572 9348
rect 12636 9284 12637 9348
rect 12571 9283 12637 9284
rect 12041 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12361 9280
rect 12041 8192 12361 9216
rect 12041 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12361 8192
rect 12041 8006 12361 8128
rect 12041 7770 12083 8006
rect 12319 7770 12361 8006
rect 11651 7580 11717 7581
rect 11651 7516 11652 7580
rect 11716 7516 11717 7580
rect 11651 7515 11717 7516
rect 11835 7580 11901 7581
rect 11835 7516 11836 7580
rect 11900 7516 11901 7580
rect 11835 7515 11901 7516
rect 12041 7104 12361 7770
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 11467 6764 11533 6765
rect 11467 6700 11468 6764
rect 11532 6700 11533 6764
rect 11467 6699 11533 6700
rect 11283 6492 11349 6493
rect 11283 6428 11284 6492
rect 11348 6428 11349 6492
rect 11283 6427 11349 6428
rect 12041 6016 12361 7040
rect 12574 6085 12634 9283
rect 12701 8736 13021 9760
rect 12701 8672 12709 8736
rect 12773 8672 12789 8736
rect 12853 8672 12869 8736
rect 12933 8672 12949 8736
rect 13013 8672 13021 8736
rect 12701 8666 13021 8672
rect 12701 8430 12743 8666
rect 12979 8430 13021 8666
rect 12701 7648 13021 8430
rect 12701 7584 12709 7648
rect 12773 7584 12789 7648
rect 12853 7584 12869 7648
rect 12933 7584 12949 7648
rect 13013 7584 13021 7648
rect 12701 6560 13021 7584
rect 12701 6496 12709 6560
rect 12773 6496 12789 6560
rect 12853 6496 12869 6560
rect 12933 6496 12949 6560
rect 13013 6496 13021 6560
rect 12571 6084 12637 6085
rect 12571 6020 12572 6084
rect 12636 6020 12637 6084
rect 12571 6019 12637 6020
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 10547 5540 10613 5541
rect 10547 5476 10548 5540
rect 10612 5476 10613 5540
rect 10547 5475 10613 5476
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 4198 12361 4864
rect 9627 4180 9693 4181
rect 9627 4116 9628 4180
rect 9692 4116 9693 4180
rect 9627 4115 9693 4116
rect 8262 3232 8270 3296
rect 8334 3232 8350 3296
rect 8414 3232 8430 3296
rect 8494 3232 8510 3296
rect 8574 3232 8582 3296
rect 8262 2208 8582 3232
rect 8262 2144 8270 2208
rect 8334 2144 8350 2208
rect 8414 2144 8430 2208
rect 8494 2144 8510 2208
rect 8574 2144 8582 2208
rect 8262 274 8582 2144
rect 8262 38 8304 274
rect 8540 38 8582 274
rect 8262 -4 8582 38
rect 12041 3962 12083 4198
rect 12319 3962 12361 4198
rect 12041 3840 12361 3962
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 934 12361 2688
rect 12041 698 12083 934
rect 12319 698 12361 934
rect 12041 -4 12361 698
rect 12701 5472 13021 6496
rect 13310 6085 13370 13771
rect 14043 13700 14109 13701
rect 14043 13636 14044 13700
rect 14108 13636 14109 13700
rect 14043 13635 14109 13636
rect 13675 11932 13741 11933
rect 13675 11868 13676 11932
rect 13740 11868 13741 11932
rect 13675 11867 13741 11868
rect 13491 9892 13557 9893
rect 13491 9828 13492 9892
rect 13556 9828 13557 9892
rect 13491 9827 13557 9828
rect 13494 7581 13554 9827
rect 13491 7580 13557 7581
rect 13491 7516 13492 7580
rect 13556 7516 13557 7580
rect 13491 7515 13557 7516
rect 13678 7037 13738 11867
rect 14046 10573 14106 13635
rect 14411 11116 14477 11117
rect 14411 11052 14412 11116
rect 14476 11052 14477 11116
rect 14411 11051 14477 11052
rect 14043 10572 14109 10573
rect 14043 10508 14044 10572
rect 14108 10508 14109 10572
rect 14043 10507 14109 10508
rect 14043 9620 14109 9621
rect 14043 9556 14044 9620
rect 14108 9556 14109 9620
rect 14043 9555 14109 9556
rect 14046 8261 14106 9555
rect 14043 8260 14109 8261
rect 14043 8196 14044 8260
rect 14108 8196 14109 8260
rect 14043 8195 14109 8196
rect 13675 7036 13741 7037
rect 13675 6972 13676 7036
rect 13740 6972 13741 7036
rect 13675 6971 13741 6972
rect 14414 6901 14474 11051
rect 14411 6900 14477 6901
rect 14411 6836 14412 6900
rect 14476 6836 14477 6900
rect 14411 6835 14477 6836
rect 13307 6084 13373 6085
rect 13307 6020 13308 6084
rect 13372 6020 13373 6084
rect 13307 6019 13373 6020
rect 14598 5949 14658 15267
rect 14782 8261 14842 15947
rect 16480 15808 16800 16832
rect 16480 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16800 15808
rect 16480 15622 16800 15744
rect 15515 15468 15581 15469
rect 15515 15404 15516 15468
rect 15580 15404 15581 15468
rect 15515 15403 15581 15404
rect 15147 13700 15213 13701
rect 15147 13636 15148 13700
rect 15212 13636 15213 13700
rect 15147 13635 15213 13636
rect 14963 11116 15029 11117
rect 14963 11052 14964 11116
rect 15028 11052 15029 11116
rect 14963 11051 15029 11052
rect 14779 8260 14845 8261
rect 14779 8196 14780 8260
rect 14844 8196 14845 8260
rect 14779 8195 14845 8196
rect 14595 5948 14661 5949
rect 14595 5884 14596 5948
rect 14660 5884 14661 5948
rect 14595 5883 14661 5884
rect 12701 5408 12709 5472
rect 12773 5408 12789 5472
rect 12853 5408 12869 5472
rect 12933 5408 12949 5472
rect 13013 5408 13021 5472
rect 12701 4858 13021 5408
rect 12701 4622 12743 4858
rect 12979 4622 13021 4858
rect 12701 4384 13021 4622
rect 12701 4320 12709 4384
rect 12773 4320 12789 4384
rect 12853 4320 12869 4384
rect 12933 4320 12949 4384
rect 13013 4320 13021 4384
rect 12701 3296 13021 4320
rect 12701 3232 12709 3296
rect 12773 3232 12789 3296
rect 12853 3232 12869 3296
rect 12933 3232 12949 3296
rect 13013 3232 13021 3296
rect 12701 2208 13021 3232
rect 14966 2957 15026 11051
rect 15150 3501 15210 13635
rect 15518 3773 15578 15403
rect 16480 15386 16522 15622
rect 16758 15386 16800 15622
rect 16480 14720 16800 15386
rect 16480 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16800 14720
rect 16480 13632 16800 14656
rect 16480 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16800 13632
rect 16480 12544 16800 13568
rect 16480 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16800 12544
rect 16480 11814 16800 12480
rect 16480 11578 16522 11814
rect 16758 11578 16800 11814
rect 16480 11456 16800 11578
rect 16480 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16800 11456
rect 16480 10368 16800 11392
rect 16480 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16800 10368
rect 16480 9280 16800 10304
rect 16480 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16800 9280
rect 16480 8192 16800 9216
rect 16990 8397 17050 18123
rect 17140 17440 17460 19310
rect 20720 19546 21040 19588
rect 20720 19310 20762 19546
rect 20998 19310 21040 19546
rect 17140 17376 17148 17440
rect 17212 17376 17228 17440
rect 17292 17376 17308 17440
rect 17372 17376 17388 17440
rect 17452 17376 17460 17440
rect 17140 16352 17460 17376
rect 20060 18886 20380 18928
rect 20060 18650 20102 18886
rect 20338 18650 20380 18886
rect 17723 17100 17789 17101
rect 17723 17036 17724 17100
rect 17788 17036 17789 17100
rect 17723 17035 17789 17036
rect 17140 16288 17148 16352
rect 17212 16288 17228 16352
rect 17292 16288 17308 16352
rect 17372 16288 17388 16352
rect 17452 16288 17460 16352
rect 17140 16282 17460 16288
rect 17140 16046 17182 16282
rect 17418 16046 17460 16282
rect 17140 15264 17460 16046
rect 17140 15200 17148 15264
rect 17212 15200 17228 15264
rect 17292 15200 17308 15264
rect 17372 15200 17388 15264
rect 17452 15200 17460 15264
rect 17140 14176 17460 15200
rect 17140 14112 17148 14176
rect 17212 14112 17228 14176
rect 17292 14112 17308 14176
rect 17372 14112 17388 14176
rect 17452 14112 17460 14176
rect 17140 13088 17460 14112
rect 17539 14108 17605 14109
rect 17539 14044 17540 14108
rect 17604 14044 17605 14108
rect 17539 14043 17605 14044
rect 17140 13024 17148 13088
rect 17212 13024 17228 13088
rect 17292 13024 17308 13088
rect 17372 13024 17388 13088
rect 17452 13024 17460 13088
rect 17140 12474 17460 13024
rect 17140 12238 17182 12474
rect 17418 12238 17460 12474
rect 17140 12000 17460 12238
rect 17140 11936 17148 12000
rect 17212 11936 17228 12000
rect 17292 11936 17308 12000
rect 17372 11936 17388 12000
rect 17452 11936 17460 12000
rect 17140 10912 17460 11936
rect 17140 10848 17148 10912
rect 17212 10848 17228 10912
rect 17292 10848 17308 10912
rect 17372 10848 17388 10912
rect 17452 10848 17460 10912
rect 17140 9824 17460 10848
rect 17140 9760 17148 9824
rect 17212 9760 17228 9824
rect 17292 9760 17308 9824
rect 17372 9760 17388 9824
rect 17452 9760 17460 9824
rect 17140 8736 17460 9760
rect 17140 8672 17148 8736
rect 17212 8672 17228 8736
rect 17292 8672 17308 8736
rect 17372 8672 17388 8736
rect 17452 8672 17460 8736
rect 17140 8666 17460 8672
rect 17140 8430 17182 8666
rect 17418 8430 17460 8666
rect 16987 8396 17053 8397
rect 16987 8332 16988 8396
rect 17052 8332 17053 8396
rect 16987 8331 17053 8332
rect 16480 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16800 8192
rect 16480 8006 16800 8128
rect 16480 7770 16522 8006
rect 16758 7770 16800 8006
rect 16480 7104 16800 7770
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 4198 16800 4864
rect 16480 3962 16522 4198
rect 16758 3962 16800 4198
rect 16480 3840 16800 3962
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 15515 3772 15581 3773
rect 15515 3708 15516 3772
rect 15580 3708 15581 3772
rect 15515 3707 15581 3708
rect 15147 3500 15213 3501
rect 15147 3436 15148 3500
rect 15212 3436 15213 3500
rect 15147 3435 15213 3436
rect 14963 2956 15029 2957
rect 14963 2892 14964 2956
rect 15028 2892 15029 2956
rect 14963 2891 15029 2892
rect 12701 2144 12709 2208
rect 12773 2144 12789 2208
rect 12853 2144 12869 2208
rect 12933 2144 12949 2208
rect 13013 2144 13021 2208
rect 12701 274 13021 2144
rect 12701 38 12743 274
rect 12979 38 13021 274
rect 12701 -4 13021 38
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 934 16800 2688
rect 16480 698 16522 934
rect 16758 698 16800 934
rect 16480 -4 16800 698
rect 17140 7648 17460 8430
rect 17140 7584 17148 7648
rect 17212 7584 17228 7648
rect 17292 7584 17308 7648
rect 17372 7584 17388 7648
rect 17452 7584 17460 7648
rect 17140 6560 17460 7584
rect 17140 6496 17148 6560
rect 17212 6496 17228 6560
rect 17292 6496 17308 6560
rect 17372 6496 17388 6560
rect 17452 6496 17460 6560
rect 17140 5472 17460 6496
rect 17542 6357 17602 14043
rect 17726 9621 17786 17035
rect 20060 15622 20380 18650
rect 20060 15386 20102 15622
rect 20338 15386 20380 15622
rect 17907 15060 17973 15061
rect 17907 14996 17908 15060
rect 17972 14996 17973 15060
rect 17907 14995 17973 14996
rect 17723 9620 17789 9621
rect 17723 9556 17724 9620
rect 17788 9556 17789 9620
rect 17723 9555 17789 9556
rect 17539 6356 17605 6357
rect 17539 6292 17540 6356
rect 17604 6292 17605 6356
rect 17539 6291 17605 6292
rect 17140 5408 17148 5472
rect 17212 5408 17228 5472
rect 17292 5408 17308 5472
rect 17372 5408 17388 5472
rect 17452 5408 17460 5472
rect 17140 4858 17460 5408
rect 17140 4622 17182 4858
rect 17418 4622 17460 4858
rect 17140 4384 17460 4622
rect 17140 4320 17148 4384
rect 17212 4320 17228 4384
rect 17292 4320 17308 4384
rect 17372 4320 17388 4384
rect 17452 4320 17460 4384
rect 17140 3296 17460 4320
rect 17140 3232 17148 3296
rect 17212 3232 17228 3296
rect 17292 3232 17308 3296
rect 17372 3232 17388 3296
rect 17452 3232 17460 3296
rect 17140 2208 17460 3232
rect 17910 3229 17970 14995
rect 20060 11814 20380 15386
rect 20060 11578 20102 11814
rect 20338 11578 20380 11814
rect 20060 8006 20380 11578
rect 20060 7770 20102 8006
rect 20338 7770 20380 8006
rect 20060 4198 20380 7770
rect 20060 3962 20102 4198
rect 20338 3962 20380 4198
rect 17907 3228 17973 3229
rect 17907 3164 17908 3228
rect 17972 3164 17973 3228
rect 17907 3163 17973 3164
rect 17140 2144 17148 2208
rect 17212 2144 17228 2208
rect 17292 2144 17308 2208
rect 17372 2144 17388 2208
rect 17452 2144 17460 2208
rect 17140 274 17460 2144
rect 20060 934 20380 3962
rect 20060 698 20102 934
rect 20338 698 20380 934
rect 20060 656 20380 698
rect 20720 16282 21040 19310
rect 20720 16046 20762 16282
rect 20998 16046 21040 16282
rect 20720 12474 21040 16046
rect 20720 12238 20762 12474
rect 20998 12238 21040 12474
rect 20720 8666 21040 12238
rect 20720 8430 20762 8666
rect 20998 8430 21040 8666
rect 20720 4858 21040 8430
rect 20720 4622 20762 4858
rect 20998 4622 21040 4858
rect 17140 38 17182 274
rect 17418 38 17460 274
rect 17140 -4 17460 38
rect 20720 274 21040 4622
rect 20720 38 20762 274
rect 20998 38 21040 274
rect 20720 -4 21040 38
<< via4 >>
rect -1034 19310 -798 19546
rect -1034 16046 -798 16282
rect -1034 12238 -798 12474
rect -1034 8430 -798 8666
rect -1034 4622 -798 4858
rect -374 18650 -138 18886
rect 3205 18650 3441 18886
rect -374 15386 -138 15622
rect -374 11578 -138 11814
rect -374 7770 -138 8006
rect -374 3962 -138 4198
rect 3865 19310 4101 19546
rect 7644 18650 7880 18886
rect 3205 15386 3441 15622
rect 3865 16046 4101 16282
rect 3205 11578 3441 11814
rect 3865 12238 4101 12474
rect 3205 7770 3441 8006
rect 3205 3962 3441 4198
rect -374 698 -138 934
rect 3205 698 3441 934
rect -1034 38 -798 274
rect 3865 8430 4101 8666
rect 3865 4622 4101 4858
rect 7644 15386 7880 15622
rect 7644 11578 7880 11814
rect 7644 7770 7880 8006
rect 7644 3962 7880 4198
rect 3865 38 4101 274
rect 7644 698 7880 934
rect 8304 19310 8540 19546
rect 8304 16046 8540 16282
rect 8304 12238 8540 12474
rect 8304 8430 8540 8666
rect 12083 18650 12319 18886
rect 8304 4622 8540 4858
rect 12083 15386 12319 15622
rect 12083 11578 12319 11814
rect 12743 19310 12979 19546
rect 12743 16046 12979 16282
rect 16522 18650 16758 18886
rect 17182 19310 17418 19546
rect 12743 12238 12979 12474
rect 12083 7770 12319 8006
rect 12743 8430 12979 8666
rect 8304 38 8540 274
rect 12083 3962 12319 4198
rect 12083 698 12319 934
rect 12743 4622 12979 4858
rect 16522 15386 16758 15622
rect 16522 11578 16758 11814
rect 20762 19310 20998 19546
rect 20102 18650 20338 18886
rect 17182 16046 17418 16282
rect 17182 12238 17418 12474
rect 17182 8430 17418 8666
rect 16522 7770 16758 8006
rect 16522 3962 16758 4198
rect 12743 38 12979 274
rect 16522 698 16758 934
rect 20102 15386 20338 15622
rect 17182 4622 17418 4858
rect 20102 11578 20338 11814
rect 20102 7770 20338 8006
rect 20102 3962 20338 4198
rect 20102 698 20338 934
rect 20762 16046 20998 16282
rect 20762 12238 20998 12474
rect 20762 8430 20998 8666
rect 20762 4622 20998 4858
rect 17182 38 17418 274
rect 20762 38 20998 274
<< metal5 >>
rect -1076 19546 21040 19588
rect -1076 19310 -1034 19546
rect -798 19310 3865 19546
rect 4101 19310 8304 19546
rect 8540 19310 12743 19546
rect 12979 19310 17182 19546
rect 17418 19310 20762 19546
rect 20998 19310 21040 19546
rect -1076 19268 21040 19310
rect -416 18886 20380 18928
rect -416 18650 -374 18886
rect -138 18650 3205 18886
rect 3441 18650 7644 18886
rect 7880 18650 12083 18886
rect 12319 18650 16522 18886
rect 16758 18650 20102 18886
rect 20338 18650 20380 18886
rect -416 18608 20380 18650
rect -1076 16282 21040 16324
rect -1076 16046 -1034 16282
rect -798 16046 3865 16282
rect 4101 16046 8304 16282
rect 8540 16046 12743 16282
rect 12979 16046 17182 16282
rect 17418 16046 20762 16282
rect 20998 16046 21040 16282
rect -1076 16004 21040 16046
rect -1076 15622 21040 15664
rect -1076 15386 -374 15622
rect -138 15386 3205 15622
rect 3441 15386 7644 15622
rect 7880 15386 12083 15622
rect 12319 15386 16522 15622
rect 16758 15386 20102 15622
rect 20338 15386 21040 15622
rect -1076 15344 21040 15386
rect -1076 12474 21040 12516
rect -1076 12238 -1034 12474
rect -798 12238 3865 12474
rect 4101 12238 8304 12474
rect 8540 12238 12743 12474
rect 12979 12238 17182 12474
rect 17418 12238 20762 12474
rect 20998 12238 21040 12474
rect -1076 12196 21040 12238
rect -1076 11814 21040 11856
rect -1076 11578 -374 11814
rect -138 11578 3205 11814
rect 3441 11578 7644 11814
rect 7880 11578 12083 11814
rect 12319 11578 16522 11814
rect 16758 11578 20102 11814
rect 20338 11578 21040 11814
rect -1076 11536 21040 11578
rect -1076 8666 21040 8708
rect -1076 8430 -1034 8666
rect -798 8430 3865 8666
rect 4101 8430 8304 8666
rect 8540 8430 12743 8666
rect 12979 8430 17182 8666
rect 17418 8430 20762 8666
rect 20998 8430 21040 8666
rect -1076 8388 21040 8430
rect -1076 8006 21040 8048
rect -1076 7770 -374 8006
rect -138 7770 3205 8006
rect 3441 7770 7644 8006
rect 7880 7770 12083 8006
rect 12319 7770 16522 8006
rect 16758 7770 20102 8006
rect 20338 7770 21040 8006
rect -1076 7728 21040 7770
rect -1076 4858 21040 4900
rect -1076 4622 -1034 4858
rect -798 4622 3865 4858
rect 4101 4622 8304 4858
rect 8540 4622 12743 4858
rect 12979 4622 17182 4858
rect 17418 4622 20762 4858
rect 20998 4622 21040 4858
rect -1076 4580 21040 4622
rect -1076 4198 21040 4240
rect -1076 3962 -374 4198
rect -138 3962 3205 4198
rect 3441 3962 7644 4198
rect 7880 3962 12083 4198
rect 12319 3962 16522 4198
rect 16758 3962 20102 4198
rect 20338 3962 21040 4198
rect -1076 3920 21040 3962
rect -416 934 20380 976
rect -416 698 -374 934
rect -138 698 3205 934
rect 3441 698 7644 934
rect 7880 698 12083 934
rect 12319 698 16522 934
rect 16758 698 20102 934
rect 20338 698 20380 934
rect -416 656 20380 698
rect -1076 274 21040 316
rect -1076 38 -1034 274
rect -798 38 3865 274
rect 4101 38 8304 274
rect 8540 38 12743 274
rect 12979 38 17182 274
rect 17418 38 20762 274
rect 20998 38 21040 274
rect -1076 -4 21040 38
use sky130_fd_sc_hd__and3_2  _151_
timestamp 0
transform -1 0 10120 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _152_
timestamp 0
transform -1 0 12696 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _153_
timestamp 0
transform 1 0 17204 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _154_
timestamp 0
transform 1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_4  _155_
timestamp 0
transform 1 0 9936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _156_
timestamp 0
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _157_
timestamp 0
transform -1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _158_
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _159_
timestamp 0
transform -1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp 0
transform -1 0 14812 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _161_
timestamp 0
transform 1 0 16192 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp 0
transform -1 0 7176 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _163_
timestamp 0
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _164_
timestamp 0
transform 1 0 4600 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _165_
timestamp 0
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 0
transform 1 0 15640 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _167_
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _168_
timestamp 0
transform -1 0 7176 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _169_
timestamp 0
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _170_
timestamp 0
transform 1 0 14444 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _171_
timestamp 0
transform -1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _172_
timestamp 0
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_4  _173_
timestamp 0
transform 1 0 6348 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _174_
timestamp 0
transform -1 0 4692 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _175_
timestamp 0
transform -1 0 7728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _176_
timestamp 0
transform -1 0 2300 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _177_
timestamp 0
transform 1 0 12512 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _178_
timestamp 0
transform -1 0 3312 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _179_
timestamp 0
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _180_
timestamp 0
transform -1 0 17572 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _181_
timestamp 0
transform 1 0 17112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _182_
timestamp 0
transform -1 0 12512 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _183_
timestamp 0
transform 1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 0
transform 1 0 2576 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _185_
timestamp 0
transform 1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 0
transform 1 0 3956 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _187_
timestamp 0
transform -1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _188_
timestamp 0
transform -1 0 10488 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _189_
timestamp 0
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_0  _190_
timestamp 0
transform -1 0 2852 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_2  _191_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _192_
timestamp 0
transform -1 0 15824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _193_
timestamp 0
transform -1 0 14996 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _194_
timestamp 0
transform -1 0 14720 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _195_
timestamp 0
transform -1 0 17112 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _196_
timestamp 0
transform -1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_4  _197_
timestamp 0
transform 1 0 8372 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _198_
timestamp 0
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_4  _199_
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_2  _200_
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_4  _201_
timestamp 0
transform -1 0 8832 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_2  _202_
timestamp 0
transform -1 0 8740 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_4  _203_
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__a22oi_4  _204_
timestamp 0
transform 1 0 16744 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_2  _205_
timestamp 0
transform -1 0 14628 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _206_
timestamp 0
transform -1 0 15548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_4  _207_
timestamp 0
transform -1 0 9108 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_2  _208_
timestamp 0
transform -1 0 7084 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _209_
timestamp 0
transform -1 0 2208 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _210_
timestamp 0
transform 1 0 16376 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__lpflow_clkinvkapwr_1  _211_
timestamp 0
transform -1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _212_
timestamp 0
transform -1 0 11960 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _213_
timestamp 0
transform -1 0 18492 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _214_
timestamp 0
transform -1 0 16100 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_8  _215_
timestamp 0
transform -1 0 3680 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_0  _216_
timestamp 0
transform -1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _217_
timestamp 0
transform -1 0 4324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _218_
timestamp 0
transform 1 0 17664 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _219_
timestamp 0
transform -1 0 7084 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _220_
timestamp 0
transform 1 0 2392 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_0  _221_
timestamp 0
transform -1 0 13156 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _222_
timestamp 0
transform -1 0 10120 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_0  _223_
timestamp 0
transform 1 0 13064 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _224_
timestamp 0
transform 1 0 15088 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _225_
timestamp 0
transform -1 0 2300 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _226_
timestamp 0
transform 1 0 8648 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _227_
timestamp 0
transform 1 0 7176 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _228_
timestamp 0
transform 1 0 11684 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_0  _229_
timestamp 0
transform -1 0 15548 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _230_
timestamp 0
transform -1 0 7176 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_0  _231_
timestamp 0
transform 1 0 13248 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _232_
timestamp 0
transform 1 0 14168 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_0  _233_
timestamp 0
transform 1 0 4140 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _234_
timestamp 0
transform 1 0 5336 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_inputiso0n_1  _235_
timestamp 0
transform -1 0 12696 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_4  _236_
timestamp 0
transform -1 0 3680 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _237_
timestamp 0
transform 1 0 1472 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_0  _238_
timestamp 0
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 0
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _240_
timestamp 0
transform 1 0 3220 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _241_
timestamp 0
transform -1 0 5888 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__or3b_4  _242_
timestamp 0
transform -1 0 2208 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _243_
timestamp 0
transform -1 0 5520 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_inputiso0n_1  _244_
timestamp 0
transform 1 0 5796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _245_
timestamp 0
transform 1 0 10856 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _246_
timestamp 0
transform 1 0 1564 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _247_
timestamp 0
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _248_
timestamp 0
transform 1 0 17756 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a2111oi_2  _249_
timestamp 0
transform 1 0 14076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ba_2  _250_
timestamp 0
transform -1 0 8556 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _251_
timestamp 0
transform 1 0 4232 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _252_
timestamp 0
transform 1 0 5888 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _253_
timestamp 0
transform 1 0 17112 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_0  _254_
timestamp 0
transform -1 0 18492 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _255_
timestamp 0
transform -1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_2  _256_
timestamp 0
transform 1 0 17572 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_inputiso0n_1  _257_
timestamp 0
transform -1 0 2392 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_clkinvkapwr_1  _258_
timestamp 0
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _259_
timestamp 0
transform 1 0 14812 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _260_
timestamp 0
transform -1 0 9200 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _261_
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _262_
timestamp 0
transform -1 0 2852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__lpflow_inputiso0n_1  _263_
timestamp 0
transform -1 0 8832 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_2  _264_
timestamp 0
transform -1 0 5152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ba_2  _265_
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__lpflow_clkinvkapwr_1  _266_
timestamp 0
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_0  _267_
timestamp 0
transform -1 0 16560 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _268_
timestamp 0
transform 1 0 11776 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _269_
timestamp 0
transform 1 0 17756 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _270_
timestamp 0
transform 1 0 17388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _271_
timestamp 0
transform 1 0 12052 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _272_
timestamp 0
transform 1 0 13984 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _273_
timestamp 0
transform 1 0 12144 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__lpflow_inputiso0n_1  _274_
timestamp 0
transform 1 0 8372 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso0n_1  _275_
timestamp 0
transform 1 0 7636 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _276_
timestamp 0
transform 1 0 4048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _277_
timestamp 0
transform 1 0 10212 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _278_
timestamp 0
transform -1 0 11408 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _279_
timestamp 0
transform -1 0 13340 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_2  _280_
timestamp 0
transform -1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ba_2  _281_
timestamp 0
transform 1 0 17848 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 0
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _283_
timestamp 0
transform -1 0 10580 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _284_
timestamp 0
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_4  _285_
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 0
transform 1 0 15364 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _287_
timestamp 0
transform 1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _288_
timestamp 0
transform -1 0 6164 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _289_
timestamp 0
transform 1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _290_
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _291_
timestamp 0
transform -1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _292_
timestamp 0
transform -1 0 7176 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _293_
timestamp 0
transform -1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _294_
timestamp 0
transform -1 0 4140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _295_
timestamp 0
transform -1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _296_
timestamp 0
transform -1 0 8004 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _297_
timestamp 0
transform 1 0 15364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _298_
timestamp 0
transform 1 0 15456 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _299_
timestamp 0
transform 1 0 14076 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _300_
timestamp 0
transform -1 0 8556 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__lpflow_clkbufkapwr_1  _301_
timestamp 0
transform 1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _302_
timestamp 0
transform 1 0 11684 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _303_
timestamp 0
transform 1 0 9292 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _304_
timestamp 0
transform 1 0 3220 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _305_
timestamp 0
transform -1 0 13432 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _306_
timestamp 0
transform 1 0 1472 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _307_
timestamp 0
transform -1 0 13616 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _308_
timestamp 0
transform 1 0 4140 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _309_
timestamp 0
transform 1 0 4140 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _310_
timestamp 0
transform 1 0 16468 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _311_
timestamp 0
transform -1 0 6348 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _312_
timestamp 0
transform -1 0 14996 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _313_
timestamp 0
transform -1 0 7636 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _314_
timestamp 0
transform -1 0 16468 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _315_
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _316_
timestamp 0
transform -1 0 16192 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _317_
timestamp 0
transform -1 0 16008 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _318_
timestamp 0
transform -1 0 3864 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _319_
timestamp 0
transform -1 0 4876 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_4  _320_
timestamp 0
transform 1 0 11776 0 -1 13056
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_2  _321_
timestamp 0
transform 1 0 7176 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _322_
timestamp 0
transform -1 0 12236 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_4  _323_
timestamp 0
transform 1 0 2944 0 -1 16320
box -38 -48 2246 592
use sky130_fd_sc_hd__dfstp_4  _324_
timestamp 0
transform 1 0 12880 0 -1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_2  _325_
timestamp 0
transform 1 0 11776 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _326_
timestamp 0
transform -1 0 6256 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _327_
timestamp 0
transform 1 0 14628 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _328_
timestamp 0
transform -1 0 3680 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _329_
timestamp 0
transform -1 0 5888 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _330_
timestamp 0
transform -1 0 11132 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _331_
timestamp 0
transform -1 0 7452 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _332_
timestamp 0
transform -1 0 8832 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _333_
timestamp 0
transform -1 0 9844 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _334_
timestamp 0
transform 1 0 11960 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _335_
timestamp 0
transform -1 0 5704 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _336_
timestamp 0
transform -1 0 10856 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_4  _337_
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_2  _338_
timestamp 0
transform 1 0 2392 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _339_
timestamp 0
transform -1 0 13524 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _340_
timestamp 0
transform 1 0 15640 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _341_
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _342_
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _343_
timestamp 0
transform -1 0 12972 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _344_
timestamp 0
transform -1 0 9476 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _345_
timestamp 0
transform 1 0 3404 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _348_
timestamp 0
transform -1 0 16468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform -1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__B
timestamp 0
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__C
timestamp 0
transform 1 0 9200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__SLEEP
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A0
timestamp 0
transform 1 0 17848 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A1
timestamp 0
transform 1 0 14996 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__S
timestamp 0
transform -1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A1
timestamp 0
transform 1 0 11132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__S
timestamp 0
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A0
timestamp 0
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A1
timestamp 0
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__S
timestamp 0
transform 1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A1
timestamp 0
transform 1 0 7360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__S
timestamp 0
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A0
timestamp 0
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A1
timestamp 0
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__S
timestamp 0
transform -1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A1
timestamp 0
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__S
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A1
timestamp 0
transform 1 0 7360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__S
timestamp 0
transform 1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A0
timestamp 0
transform -1 0 13984 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A1
timestamp 0
transform -1 0 14444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__S
timestamp 0
transform -1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A
timestamp 0
transform -1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A0
timestamp 0
transform 1 0 5336 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A1
timestamp 0
transform 1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__S
timestamp 0
transform 1 0 6440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A0
timestamp 0
transform -1 0 2668 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A1
timestamp 0
transform 1 0 2668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__S
timestamp 0
transform 1 0 2852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A0
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A1
timestamp 0
transform 1 0 4416 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__S
timestamp 0
transform -1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A1
timestamp 0
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__S
timestamp 0
transform 1 0 16560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A1
timestamp 0
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__S
timestamp 0
transform 1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A0
timestamp 0
transform -1 0 2944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A1
timestamp 0
transform -1 0 3680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__S
timestamp 0
transform 1 0 2392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A1
timestamp 0
transform -1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__S
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A1
timestamp 0
transform 1 0 9108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__S
timestamp 0
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 0
transform -1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A1
timestamp 0
transform -1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A2
timestamp 0
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 0
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A2
timestamp 0
transform -1 0 14720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B1_N
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A1
timestamp 0
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A2
timestamp 0
transform -1 0 13892 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 0
transform -1 0 17848 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__B
timestamp 0
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 0
transform 1 0 6164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__B
timestamp 0
transform 1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__C
timestamp 0
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A1
timestamp 0
transform 1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A2
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__B2
timestamp 0
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A1
timestamp 0
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A2
timestamp 0
transform 1 0 12696 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__B1
timestamp 0
transform 1 0 12696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__B2
timestamp 0
transform 1 0 15180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 0
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__B
timestamp 0
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__C
timestamp 0
transform 1 0 11592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__D
timestamp 0
transform 1 0 11224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A1
timestamp 0
transform 1 0 7820 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A2
timestamp 0
transform -1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__B1
timestamp 0
transform -1 0 9292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__B2
timestamp 0
transform 1 0 7820 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 0
transform 1 0 5520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__B
timestamp 0
transform 1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__C
timestamp 0
transform 1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__D
timestamp 0
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A1
timestamp 0
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A2
timestamp 0
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__B1
timestamp 0
transform 1 0 16008 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__B2
timestamp 0
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 0
transform -1 0 15180 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__B
timestamp 0
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__C
timestamp 0
transform -1 0 14444 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__D
timestamp 0
transform -1 0 13984 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__C1
timestamp 0
transform -1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A2
timestamp 0
transform 1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A2
timestamp 0
transform -1 0 7268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__B1
timestamp 0
transform -1 0 8004 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__C1
timestamp 0
transform -1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 0
transform 1 0 2944 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__B
timestamp 0
transform 1 0 3036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__C
timestamp 0
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__D
timestamp 0
transform 1 0 2576 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 0
transform 1 0 16008 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__B
timestamp 0
transform 1 0 16192 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__C
timestamp 0
transform -1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__D
timestamp 0
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 0
transform -1 0 9476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A1
timestamp 0
transform -1 0 17756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A2
timestamp 0
transform -1 0 17388 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__C1
timestamp 0
transform 1 0 17572 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__B
timestamp 0
transform -1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 0
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__B
timestamp 0
transform 1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A1
timestamp 0
transform -1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A2
timestamp 0
transform 1 0 17204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__B1
timestamp 0
transform -1 0 17480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A1
timestamp 0
transform 1 0 7912 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A2
timestamp 0
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__B1
timestamp 0
transform 1 0 7268 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__B2
timestamp 0
transform 1 0 8280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 0
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__B
timestamp 0
transform -1 0 3588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 0
transform 1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__B
timestamp 0
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1
timestamp 0
transform 1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B1
timestamp 0
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B2
timestamp 0
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 0
transform 1 0 12788 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__B
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A1
timestamp 0
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A2
timestamp 0
transform 1 0 14076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__B1
timestamp 0
transform -1 0 17204 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__B2
timestamp 0
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 0
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__B
timestamp 0
transform -1 0 2392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__C
timestamp 0
transform 1 0 2852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A1
timestamp 0
transform 1 0 8464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__B1
timestamp 0
transform 1 0 8280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__B2
timestamp 0
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 0
transform 1 0 6992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__B
timestamp 0
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__C
timestamp 0
transform -1 0 8096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A1
timestamp 0
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A2
timestamp 0
transform -1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__B1
timestamp 0
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__B2
timestamp 0
transform -1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 0
transform 1 0 14720 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__B
timestamp 0
transform 1 0 16652 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A1
timestamp 0
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__B1
timestamp 0
transform 1 0 5336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__B2
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 0
transform 1 0 12880 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B
timestamp 0
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A1
timestamp 0
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__B1
timestamp 0
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__B2
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 0
transform -1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__B
timestamp 0
transform -1 0 3680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 0
transform 1 0 5152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A2
timestamp 0
transform 1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B1
timestamp 0
transform -1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B2
timestamp 0
transform 1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 0
transform 1 0 13248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__SLEEP_B
timestamp 0
transform 1 0 12880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 0
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A2
timestamp 0
transform 1 0 2208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 0
transform -1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__SLEEP
timestamp 0
transform -1 0 6256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 0
transform 1 0 4508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__SLEEP_B
timestamp 0
transform 1 0 5244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 0
transform 1 0 10672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 0
transform 1 0 3404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__B
timestamp 0
transform -1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A1
timestamp 0
transform -1 0 6716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A2
timestamp 0
transform -1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B1
timestamp 0
transform -1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B2
timestamp 0
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 0
transform -1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__B
timestamp 0
transform -1 0 17756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A1
timestamp 0
transform 1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A2
timestamp 0
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__D1
timestamp 0
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A2
timestamp 0
transform -1 0 7636 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__D_N
timestamp 0
transform 1 0 4048 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__SLEEP
timestamp 0
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 0
transform 1 0 16744 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__B
timestamp 0
transform 1 0 16928 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A1
timestamp 0
transform 1 0 17940 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__B1
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A1
timestamp 0
transform -1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A2
timestamp 0
transform -1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__B1
timestamp 0
transform -1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A3
timestamp 0
transform -1 0 15824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__B1
timestamp 0
transform 1 0 18124 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__B2
timestamp 0
transform 1 0 17020 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 0
transform -1 0 2760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__SLEEP_B
timestamp 0
transform 1 0 2392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 0
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A2
timestamp 0
transform 1 0 14628 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__B1
timestamp 0
transform 1 0 14628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A1
timestamp 0
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A2
timestamp 0
transform 1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__B1
timestamp 0
transform 1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__B2
timestamp 0
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A2
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A1
timestamp 0
transform 1 0 3220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A2
timestamp 0
transform 1 0 2852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__B1
timestamp 0
transform 1 0 3036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 0
transform -1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__SLEEP_B
timestamp 0
transform -1 0 8372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A2
timestamp 0
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__D1
timestamp 0
transform 1 0 5336 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A1
timestamp 0
transform 1 0 16008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A2
timestamp 0
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__B1
timestamp 0
transform 1 0 17296 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A
timestamp 0
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__SLEEP
timestamp 0
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A1
timestamp 0
transform 1 0 17296 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A2
timestamp 0
transform -1 0 17572 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__B1
timestamp 0
transform -1 0 17940 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__B2
timestamp 0
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A1
timestamp 0
transform -1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A2
timestamp 0
transform 1 0 17572 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A1
timestamp 0
transform -1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A2
timestamp 0
transform -1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__B1
timestamp 0
transform -1 0 12052 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__B2
timestamp 0
transform -1 0 13524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A2
timestamp 0
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__B1
timestamp 0
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__B2
timestamp 0
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__C1
timestamp 0
transform 1 0 14444 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A1
timestamp 0
transform 1 0 12880 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A2
timestamp 0
transform 1 0 11960 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__SLEEP_B
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 0
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__SLEEP_B
timestamp 0
transform 1 0 8096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A1
timestamp 0
transform 1 0 5244 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A2
timestamp 0
transform 1 0 5980 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__B1
timestamp 0
transform 1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__C1
timestamp 0
transform 1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__B1
timestamp 0
transform -1 0 10212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__B2
timestamp 0
transform 1 0 9844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A1
timestamp 0
transform 1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A2
timestamp 0
transform 1 0 10488 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__B1
timestamp 0
transform 1 0 10120 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__B2
timestamp 0
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 0
transform 1 0 12512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__SLEEP
timestamp 0
transform 1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A2
timestamp 0
transform 1 0 6716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__D1
timestamp 0
transform -1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A1
timestamp 0
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A2
timestamp 0
transform 1 0 17664 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A
timestamp 0
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A2
timestamp 0
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__B
timestamp 0
transform -1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A0
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A1
timestamp 0
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__S
timestamp 0
transform 1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A1
timestamp 0
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__S
timestamp 0
transform -1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 0
transform 1 0 16836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A0
timestamp 0
transform 1 0 4600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A1
timestamp 0
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__S
timestamp 0
transform 1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A0
timestamp 0
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A1
timestamp 0
transform 1 0 7728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__S
timestamp 0
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A0
timestamp 0
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A1
timestamp 0
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__S
timestamp 0
transform 1 0 4048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A0
timestamp 0
transform 1 0 8740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A1
timestamp 0
transform 1 0 8372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__S
timestamp 0
transform 1 0 8556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A0
timestamp 0
transform 1 0 15548 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A1
timestamp 0
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__S
timestamp 0
transform 1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A0
timestamp 0
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A1
timestamp 0
transform -1 0 7544 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__S
timestamp 0
transform -1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__SET_B
timestamp 0
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__D
timestamp 0
transform 1 0 5336 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__RESET_B
timestamp 0
transform 1 0 14536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__D
timestamp 0
transform -1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__RESET_B
timestamp 0
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__D
timestamp 0
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__D
timestamp 0
transform -1 0 5060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__SET_B
timestamp 0
transform 1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__SET_B
timestamp 0
transform -1 0 15824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__D
timestamp 0
transform -1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__RESET_B
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__RESET_B
timestamp 0
transform 1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__D
timestamp 0
transform 1 0 5704 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__SET_B
timestamp 0
transform -1 0 16284 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__RESET_B
timestamp 0
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__D
timestamp 0
transform -1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__RESET_B
timestamp 0
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__SET_B
timestamp 0
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 0
transform -1 0 16560 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 0
transform 1 0 9292 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout38_A
timestamp 0
transform 1 0 6072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout39_A
timestamp 0
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout40_A
timestamp 0
transform 1 0 12972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 0
transform -1 0 2300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 0
transform -1 0 4508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 0
transform -1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 0
transform -1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 0
transform -1 0 3404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 0
transform -1 0 3220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 0
transform -1 0 2392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 0
transform -1 0 2944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 0
transform -1 0 2576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 0
transform -1 0 2024 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 0
transform -1 0 3864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 0
transform -1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 0
transform -1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 0
transform -1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 0
transform -1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 0
transform -1 0 12328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 0
transform -1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 0
transform -1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 0
transform -1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 0
transform -1 0 8556 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 0
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 0
transform -1 0 11408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output23_A
timestamp 0
transform 1 0 5704 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output24_A
timestamp 0
transform -1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output25_A
timestamp 0
transform 1 0 2668 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_A
timestamp 0
transform -1 0 2576 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output29_A
timestamp 0
transform -1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 0
transform -1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 0
transform -1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output32_A
timestamp 0
transform 1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output33_A
timestamp 0
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 9476 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 8188 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform -1 0 7820 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform 1 0 12144 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 12788 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinvlp_4  clkload0
timestamp 0
transform 1 0 6256 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  clkload1
timestamp 0
transform 1 0 5704 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 0
transform 1 0 12788 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout36
timestamp 0
transform -1 0 2944 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout37
timestamp 0
transform 1 0 4692 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 0
transform -1 0 6072 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout39
timestamp 0
transform -1 0 11040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout40
timestamp 0
transform -1 0 13340 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_17
timestamp 0
transform 1 0 2668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 0
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_33
timestamp 0
transform 1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_61
timestamp 0
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_65
timestamp 0
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_91
timestamp 0
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_98
timestamp 0
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_105
timestamp 0
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_144
timestamp 0
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_148
timestamp 0
transform 1 0 14720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_157
timestamp 0
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_161
timestamp 0
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 0
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_175
timestamp 0
transform 1 0 17204 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_178
timestamp 0
transform 1 0 17480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_182
timestamp 0
transform 1 0 17848 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_12
timestamp 0
transform 1 0 2208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_19
timestamp 0
transform 1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_23
timestamp 0
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_35
timestamp 0
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_43
timestamp 0
transform 1 0 5060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_46
timestamp 0
transform 1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_50
timestamp 0
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_65
timestamp 0
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_87
timestamp 0
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_91
timestamp 0
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_95
timestamp 0
transform 1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_108
timestamp 0
transform 1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_121
timestamp 0
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_152
timestamp 0
transform 1 0 15088 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_156
timestamp 0
transform 1 0 15456 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_160
timestamp 0
transform 1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 0
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_173
timestamp 0
transform 1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_177
timestamp 0
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_187
timestamp 0
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_9
timestamp 0
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_13
timestamp 0
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_18
timestamp 0
transform 1 0 2760 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_22
timestamp 0
transform 1 0 3128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_38
timestamp 0
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_43
timestamp 0
transform 1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_55
timestamp 0
transform 1 0 6164 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_59
timestamp 0
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_71
timestamp 0
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_76
timestamp 0
transform 1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 0
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_89
timestamp 0
transform 1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_93
timestamp 0
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_117
timestamp 0
transform 1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_122
timestamp 0
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_128
timestamp 0
transform 1 0 12880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_138
timestamp 0
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_151
timestamp 0
transform 1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_155
timestamp 0
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_11
timestamp 0
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_52
timestamp 0
transform 1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_87
timestamp 0
transform 1 0 9108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 0
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_151
timestamp 0
transform 1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_155
timestamp 0
transform 1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_159
timestamp 0
transform 1 0 15732 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_165
timestamp 0
transform 1 0 16284 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_9
timestamp 0
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_13
timestamp 0
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_17
timestamp 0
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_23
timestamp 0
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_51
timestamp 0
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_55
timestamp 0
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_67
timestamp 0
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_137
timestamp 0
transform 1 0 13708 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_144
timestamp 0
transform 1 0 14352 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_148
timestamp 0
transform 1 0 14720 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_160
timestamp 0
transform 1 0 15824 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_168
timestamp 0
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_176
timestamp 0
transform 1 0 17296 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_185
timestamp 0
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_189
timestamp 0
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_9
timestamp 0
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_44
timestamp 0
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 0
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_61
timestamp 0
transform 1 0 6716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_67
timestamp 0
transform 1 0 7268 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_70
timestamp 0
transform 1 0 7544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_95
timestamp 0
transform 1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_100
timestamp 0
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_183
timestamp 0
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_189
timestamp 0
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_13
timestamp 0
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_18
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_22
timestamp 0
transform 1 0 3128 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_33
timestamp 0
transform 1 0 4140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_45
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_48
timestamp 0
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_66
timestamp 0
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_70
timestamp 0
transform 1 0 7544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_74
timestamp 0
transform 1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_79
timestamp 0
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_91
timestamp 0
transform 1 0 9476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_103
timestamp 0
transform 1 0 10580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_115
timestamp 0
transform 1 0 11684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_123
timestamp 0
transform 1 0 12420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_126
timestamp 0
transform 1 0 12696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_130
timestamp 0
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 0
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_162
timestamp 0
transform 1 0 16008 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_174
timestamp 0
transform 1 0 17112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_178
timestamp 0
transform 1 0 17480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_181
timestamp 0
transform 1 0 17756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_185
timestamp 0
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_9
timestamp 0
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_24
timestamp 0
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_30
timestamp 0
transform 1 0 3864 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_34
timestamp 0
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_38
timestamp 0
transform 1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_42
timestamp 0
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 0
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_66
timestamp 0
transform 1 0 7176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_94
timestamp 0
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_102
timestamp 0
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 0
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 0
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_133
timestamp 0
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_175
timestamp 0
transform 1 0 17204 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_179
timestamp 0
transform 1 0 17572 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_183
timestamp 0
transform 1 0 17940 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_187
timestamp 0
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_12
timestamp 0
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_21
timestamp 0
transform 1 0 3036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_38
timestamp 0
transform 1 0 4600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_69
timestamp 0
transform 1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_93
timestamp 0
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_96
timestamp 0
transform 1 0 9936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_131
timestamp 0
transform 1 0 13156 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_135
timestamp 0
transform 1 0 13524 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_145
timestamp 0
transform 1 0 14444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_157
timestamp 0
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_170
timestamp 0
transform 1 0 16744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_174
timestamp 0
transform 1 0 17112 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_178
timestamp 0
transform 1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_30
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_34
timestamp 0
transform 1 0 4232 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_48
timestamp 0
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_87
timestamp 0
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_90
timestamp 0
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_94
timestamp 0
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_106
timestamp 0
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 0
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_119
timestamp 0
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_149
timestamp 0
transform 1 0 14812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_153
timestamp 0
transform 1 0 15180 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_156
timestamp 0
transform 1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_160
timestamp 0
transform 1 0 15824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_164
timestamp 0
transform 1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_188
timestamp 0
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_19
timestamp 0
transform 1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_23
timestamp 0
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_46
timestamp 0
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_50
timestamp 0
transform 1 0 5704 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_54
timestamp 0
transform 1 0 6072 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_58
timestamp 0
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_70
timestamp 0
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_98
timestamp 0
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_108
timestamp 0
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_112
timestamp 0
transform 1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_116
timestamp 0
transform 1 0 11776 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_128
timestamp 0
transform 1 0 12880 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_136
timestamp 0
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_145
timestamp 0
transform 1 0 14444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_163
timestamp 0
transform 1 0 16100 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_167
timestamp 0
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_172
timestamp 0
transform 1 0 16928 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_177
timestamp 0
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_181
timestamp 0
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_187
timestamp 0
transform 1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_12
timestamp 0
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_16
timestamp 0
transform 1 0 2576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_28
timestamp 0
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 0
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_77
timestamp 0
transform 1 0 8188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_87
timestamp 0
transform 1 0 9108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_134
timestamp 0
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_138
timestamp 0
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_142
timestamp 0
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_146
timestamp 0
transform 1 0 14536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_149
timestamp 0
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_153
timestamp 0
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_164
timestamp 0
transform 1 0 16192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_179
timestamp 0
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_6
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_17
timestamp 0
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 0
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_40
timestamp 0
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_44
timestamp 0
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_47
timestamp 0
transform 1 0 5428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_62
timestamp 0
transform 1 0 6808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_102
timestamp 0
transform 1 0 10488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 0
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_144
timestamp 0
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_148
timestamp 0
transform 1 0 14720 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_152
timestamp 0
transform 1 0 15088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_155
timestamp 0
transform 1 0 15364 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_160
timestamp 0
transform 1 0 15824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_188
timestamp 0
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_26
timestamp 0
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_30
timestamp 0
transform 1 0 3864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_34
timestamp 0
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_38
timestamp 0
transform 1 0 4600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_41
timestamp 0
transform 1 0 4876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_45
timestamp 0
transform 1 0 5244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 0
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_65
timestamp 0
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_87
timestamp 0
transform 1 0 9108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_92
timestamp 0
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_96
timestamp 0
transform 1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_100
timestamp 0
transform 1 0 10304 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_139
timestamp 0
transform 1 0 13892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_153
timestamp 0
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_157
timestamp 0
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_161
timestamp 0
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 0
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_185
timestamp 0
transform 1 0 18124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 0
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_12
timestamp 0
transform 1 0 2208 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_20
timestamp 0
transform 1 0 2944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_24
timestamp 0
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_57
timestamp 0
transform 1 0 6348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_61
timestamp 0
transform 1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_72
timestamp 0
transform 1 0 7728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_76
timestamp 0
transform 1 0 8096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_79
timestamp 0
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_118
timestamp 0
transform 1 0 11960 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_126
timestamp 0
transform 1 0 12696 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_130
timestamp 0
transform 1 0 13064 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_134
timestamp 0
transform 1 0 13432 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_167
timestamp 0
transform 1 0 16468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_187
timestamp 0
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_13
timestamp 0
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_17
timestamp 0
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_21
timestamp 0
transform 1 0 3036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_71
timestamp 0
transform 1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_75
timestamp 0
transform 1 0 8004 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_78
timestamp 0
transform 1 0 8280 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_96
timestamp 0
transform 1 0 9936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_100
timestamp 0
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_104
timestamp 0
transform 1 0 10672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_108
timestamp 0
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_122
timestamp 0
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_126
timestamp 0
transform 1 0 12696 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_147
timestamp 0
transform 1 0 14628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_151
timestamp 0
transform 1 0 14996 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_159
timestamp 0
transform 1 0 15732 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_164
timestamp 0
transform 1 0 16192 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_173
timestamp 0
transform 1 0 17020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_177
timestamp 0
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_180
timestamp 0
transform 1 0 17664 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_6
timestamp 0
transform 1 0 1656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_33
timestamp 0
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_36
timestamp 0
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_40
timestamp 0
transform 1 0 4784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_44
timestamp 0
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_48
timestamp 0
transform 1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_79
timestamp 0
transform 1 0 8372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_89
timestamp 0
transform 1 0 9292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_101
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_113
timestamp 0
transform 1 0 11500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_125
timestamp 0
transform 1 0 12604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 0
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_151
timestamp 0
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_155
timestamp 0
transform 1 0 15364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_159
timestamp 0
transform 1 0 15732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_163
timestamp 0
transform 1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_173
timestamp 0
transform 1 0 17020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_182
timestamp 0
transform 1 0 17848 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_19
timestamp 0
transform 1 0 2852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_25
timestamp 0
transform 1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_36
timestamp 0
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_42
timestamp 0
transform 1 0 4968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_48
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_52
timestamp 0
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_75
timestamp 0
transform 1 0 8004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_85
timestamp 0
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_97
timestamp 0
transform 1 0 10028 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_103
timestamp 0
transform 1 0 10580 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_106
timestamp 0
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_130
timestamp 0
transform 1 0 13064 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_174
timestamp 0
transform 1 0 17112 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_178
timestamp 0
transform 1 0 17480 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_182
timestamp 0
transform 1 0 17848 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_14
timestamp 0
transform 1 0 2392 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_18
timestamp 0
transform 1 0 2760 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_23
timestamp 0
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_44
timestamp 0
transform 1 0 5152 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_48
timestamp 0
transform 1 0 5520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_117
timestamp 0
transform 1 0 11868 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_129
timestamp 0
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_136
timestamp 0
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_145
timestamp 0
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_149
timestamp 0
transform 1 0 14812 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_156
timestamp 0
transform 1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_179
timestamp 0
transform 1 0 17572 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_187
timestamp 0
transform 1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_61
timestamp 0
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_65
timestamp 0
transform 1 0 7084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_71
timestamp 0
transform 1 0 7636 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_83
timestamp 0
transform 1 0 8740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_89
timestamp 0
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_102
timestamp 0
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 0
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_149
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 0
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_180
timestamp 0
transform 1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_184
timestamp 0
transform 1 0 18032 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_12
timestamp 0
transform 1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_16
timestamp 0
transform 1 0 2576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_35
timestamp 0
transform 1 0 4324 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_57
timestamp 0
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_69
timestamp 0
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_75
timestamp 0
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_89
timestamp 0
transform 1 0 9292 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_93
timestamp 0
transform 1 0 9660 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_105
timestamp 0
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_111
timestamp 0
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_124
timestamp 0
transform 1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_128
timestamp 0
transform 1 0 12880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_134
timestamp 0
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 0
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_145
timestamp 0
transform 1 0 14444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_150
timestamp 0
transform 1 0 14904 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_161
timestamp 0
transform 1 0 15916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_167
timestamp 0
transform 1 0 16468 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_171
timestamp 0
transform 1 0 16836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_175
timestamp 0
transform 1 0 17204 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_179
timestamp 0
transform 1 0 17572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_187
timestamp 0
transform 1 0 18308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_6
timestamp 0
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_11
timestamp 0
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_16
timestamp 0
transform 1 0 2576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_20
timestamp 0
transform 1 0 2944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_41
timestamp 0
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_47
timestamp 0
transform 1 0 5428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_63
timestamp 0
transform 1 0 6900 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_66
timestamp 0
transform 1 0 7176 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_74
timestamp 0
transform 1 0 7912 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_82
timestamp 0
transform 1 0 8648 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_85
timestamp 0
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_98
timestamp 0
transform 1 0 10120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_102
timestamp 0
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 0
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_117
timestamp 0
transform 1 0 11868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_129
timestamp 0
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_135
timestamp 0
transform 1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_139
timestamp 0
transform 1 0 13892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_143
timestamp 0
transform 1 0 14260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_173
timestamp 0
transform 1 0 17020 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_185
timestamp 0
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 0
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_6
timestamp 0
transform 1 0 1656 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_10
timestamp 0
transform 1 0 2024 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_14
timestamp 0
transform 1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_19
timestamp 0
transform 1 0 2852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_23
timestamp 0
transform 1 0 3220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_54
timestamp 0
transform 1 0 6072 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_63
timestamp 0
transform 1 0 6900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_72
timestamp 0
transform 1 0 7728 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_76
timestamp 0
transform 1 0 8096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_80
timestamp 0
transform 1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_106
timestamp 0
transform 1 0 10856 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_135
timestamp 0
transform 1 0 13524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_148
timestamp 0
transform 1 0 14720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_167
timestamp 0
transform 1 0 16468 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_179
timestamp 0
transform 1 0 17572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_187
timestamp 0
transform 1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_13
timestamp 0
transform 1 0 2300 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_35
timestamp 0
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_65
timestamp 0
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_78
timestamp 0
transform 1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_91
timestamp 0
transform 1 0 9476 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_103
timestamp 0
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_117
timestamp 0
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_147
timestamp 0
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_151
timestamp 0
transform 1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_155
timestamp 0
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_159
timestamp 0
transform 1 0 15732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_163
timestamp 0
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_177
timestamp 0
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_189
timestamp 0
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_7
timestamp 0
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_13
timestamp 0
transform 1 0 2300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_17
timestamp 0
transform 1 0 2668 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_21
timestamp 0
transform 1 0 3036 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_25
timestamp 0
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_33
timestamp 0
transform 1 0 4140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_37
timestamp 0
transform 1 0 4508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_45
timestamp 0
transform 1 0 5244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_57
timestamp 0
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_63
timestamp 0
transform 1 0 6900 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_67
timestamp 0
transform 1 0 7268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_71
timestamp 0
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_75
timestamp 0
transform 1 0 8004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_80
timestamp 0
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_136
timestamp 0
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_145
timestamp 0
transform 1 0 14444 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_149
timestamp 0
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_173
timestamp 0
transform 1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_189
timestamp 0
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_9
timestamp 0
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_13
timestamp 0
transform 1 0 2300 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_16
timestamp 0
transform 1 0 2576 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_44
timestamp 0
transform 1 0 5152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_48
timestamp 0
transform 1 0 5520 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_52
timestamp 0
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_66
timestamp 0
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_70
timestamp 0
transform 1 0 7544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_75
timestamp 0
transform 1 0 8004 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_88
timestamp 0
transform 1 0 9200 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_92
timestamp 0
transform 1 0 9568 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_96
timestamp 0
transform 1 0 9936 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_108
timestamp 0
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_133
timestamp 0
transform 1 0 13340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_138
timestamp 0
transform 1 0 13800 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_144
timestamp 0
transform 1 0 14352 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_152
timestamp 0
transform 1 0 15088 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_160
timestamp 0
transform 1 0 15824 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 0
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_189
timestamp 0
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_14
timestamp 0
transform 1 0 2392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_45
timestamp 0
transform 1 0 5244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_49
timestamp 0
transform 1 0 5612 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_52
timestamp 0
transform 1 0 5888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_56
timestamp 0
transform 1 0 6256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_60
timestamp 0
transform 1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_64
timestamp 0
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_68
timestamp 0
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_72
timestamp 0
transform 1 0 7728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_75
timestamp 0
transform 1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_93
timestamp 0
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_101
timestamp 0
transform 1 0 10396 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_111
timestamp 0
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_115
timestamp 0
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_127
timestamp 0
transform 1 0 12788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_131
timestamp 0
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_135
timestamp 0
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_154
timestamp 0
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_160
timestamp 0
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_164
timestamp 0
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_173
timestamp 0
transform 1 0 17020 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_185
timestamp 0
transform 1 0 18124 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_189
timestamp 0
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_22
timestamp 0
transform 1 0 3128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 0
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_65
timestamp 0
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_72
timestamp 0
transform 1 0 7728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_76
timestamp 0
transform 1 0 8096 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_80
timestamp 0
transform 1 0 8464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_85
timestamp 0
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_89
timestamp 0
transform 1 0 9292 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_101
timestamp 0
transform 1 0 10396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_109
timestamp 0
transform 1 0 11132 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_121
timestamp 0
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_129
timestamp 0
transform 1 0 12972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_135
timestamp 0
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_139
timestamp 0
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_141
timestamp 0
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_145
timestamp 0
transform 1 0 14444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_157
timestamp 0
transform 1 0 15548 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_163
timestamp 0
transform 1 0 16100 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 0
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_189
timestamp 0
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 0
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform -1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform -1 0 2852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform -1 0 3128 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform 1 0 1932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 0
transform -1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 0
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 0
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 0
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 0
transform -1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 0
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  lfsr_axi_top_41
timestamp 0
transform -1 0 2208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  lfsr_axi_top_42
timestamp 0
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 0
transform -1 0 1932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 0
transform -1 0 1932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 0
transform -1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 0
transform -1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 0
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output28
timestamp 0
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output29
timestamp 0
transform -1 0 1932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output30
timestamp 0
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output31
timestamp 0
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output32
timestamp 0
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output33
timestamp 0
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output34
timestamp 0
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output35
timestamp 0
transform -1 0 12236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_69
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_89
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_92
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_93
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_95
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_96
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_98
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_99
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_101
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_102
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_104
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_105
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_107
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_108
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_110
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_111
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_113
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_114
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_116
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_117
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_119
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_120
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_122
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_123
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_125
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_126
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_128
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_129
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_131
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_132
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_134
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_135
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_137
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_138
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_140
timestamp 0
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_141
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 0
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 0
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
<< labels >>
rlabel metal1 s 9982 17408 9982 17408 4 VGND
rlabel metal1 s 9982 16864 9982 16864 4 VPWR
rlabel metal2 s 9108 13940 9108 13940 4 _000_
rlabel metal2 s 4462 4352 4462 4352 4 _001_
rlabel metal1 s 17434 13430 17434 13430 4 _002_
rlabel metal2 s 12650 7956 12650 7956 4 _003_
rlabel metal2 s 2254 15691 2254 15691 4 _004_
rlabel metal1 s 13754 2278 13754 2278 4 _005_
rlabel metal2 s 5198 9197 5198 9197 4 _006_
rlabel metal1 s 1840 3978 1840 3978 4 _007_
rlabel metal3 s 8234 10013 8234 10013 4 _008_
rlabel metal2 s 12558 15759 12558 15759 4 _009_
rlabel metal1 s 14490 4046 14490 4046 4 _010_
rlabel metal2 s 16836 10132 16836 10132 4 _011_
rlabel metal1 s 16514 9962 16514 9962 4 _012_
rlabel metal1 s 1748 13158 1748 13158 4 _013_
rlabel metal1 s 14582 12070 14582 12070 4 _014_
rlabel metal2 s 13938 7548 13938 7548 4 _015_
rlabel metal3 s 690 16660 690 16660 4 _016_
rlabel metal1 s 14490 14586 14490 14586 4 _017_
rlabel metal2 s 12190 12852 12190 12852 4 _018_
rlabel metal1 s 9016 13838 9016 13838 4 _019_
rlabel metal1 s 15364 13158 15364 13158 4 _020_
rlabel metal1 s 9292 15130 9292 15130 4 _021_
rlabel metal3 s 13593 7004 13593 7004 4 _022_
rlabel metal2 s 12098 2108 12098 2108 4 _023_
rlabel metal1 s 5014 2482 5014 2482 4 _024_
rlabel metal2 s 14950 13753 14950 13753 4 _025_
rlabel metal1 s 2576 9146 2576 9146 4 _026_
rlabel metal1 s 7130 8398 7130 8398 4 _027_
rlabel metal2 s 12650 4930 12650 4930 4 _028_
rlabel metal2 s 2622 8432 2622 8432 4 _029_
rlabel metal2 s 10718 9078 10718 9078 4 _030_
rlabel metal2 s 15686 7089 15686 7089 4 _031_
rlabel metal1 s 11868 15062 11868 15062 4 _032_
rlabel metal2 s 5842 16711 5842 16711 4 _033_
rlabel metal1 s 17434 10778 17434 10778 4 _034_
rlabel metal1 s 16468 3502 16468 3502 4 _035_
rlabel metal3 s 1771 14076 1771 14076 4 _036_
rlabel metal1 s 17618 14382 17618 14382 4 _037_
rlabel metal3 s 15962 12291 15962 12291 4 _038_
rlabel metal1 s 16744 4114 16744 4114 4 _039_
rlabel metal2 s 9338 15351 9338 15351 4 _040_
rlabel metal1 s 12604 8942 12604 8942 4 _041_
rlabel metal1 s 13340 16218 13340 16218 4 _042_
rlabel metal2 s 1058 8653 1058 8653 4 _043_
rlabel metal1 s 3450 2958 3450 2958 4 _044_
rlabel metal1 s 7222 10438 7222 10438 4 _045_
rlabel metal1 s 6992 10778 6992 10778 4 _046_
rlabel metal2 s 10074 8398 10074 8398 4 _047_
rlabel metal2 s 12466 16864 12466 16864 4 _048_
rlabel metal2 s 8510 12427 8510 12427 4 _049_
rlabel metal2 s 4278 4964 4278 4964 4 _050_
rlabel metal1 s 15134 7514 15134 7514 4 _051_
rlabel metal1 s 8878 16218 8878 16218 4 _052_
rlabel metal4 s 2668 10880 2668 10880 4 _053_
rlabel metal1 s 18032 2346 18032 2346 4 _054_
rlabel metal2 s 7130 7191 7130 7191 4 _055_
rlabel metal4 s 14605 15300 14605 15300 4 _056_
rlabel metal2 s 6486 14586 6486 14586 4 _057_
rlabel metal1 s 2714 6188 2714 6188 4 _058_
rlabel metal1 s 7452 10030 7452 10030 4 _059_
rlabel metal3 s 12742 16099 12742 16099 4 _060_
rlabel metal1 s 4232 6426 4232 6426 4 _061_
rlabel metal2 s 17526 7684 17526 7684 4 _062_
rlabel metal1 s 16514 16014 16514 16014 4 _063_
rlabel metal2 s 1886 14858 1886 14858 4 _064_
rlabel metal2 s 3082 6154 3082 6154 4 _065_
rlabel metal2 s 13616 10948 13616 10948 4 _066_
rlabel metal2 s 3174 3026 3174 3026 4 _067_
rlabel metal2 s 15410 17119 15410 17119 4 _068_
rlabel metal4 s 14421 11084 14421 11084 4 _069_
rlabel metal1 s 2300 10438 2300 10438 4 _070_
rlabel metal3 s 15042 9724 15042 9724 4 _071_
rlabel metal3 s 12604 10812 12604 10812 4 _072_
rlabel metal2 s 13662 4114 13662 4114 4 _073_
rlabel metal1 s 9246 4658 9246 4658 4 _074_
rlabel metal2 s 17894 15181 17894 15181 4 _075_
rlabel metal2 s 17526 5389 17526 5389 4 _076_
rlabel metal2 s 15134 2244 15134 2244 4 _077_
rlabel metal1 s 9200 2482 9200 2482 4 _078_
rlabel metal1 s 11914 2584 11914 2584 4 _079_
rlabel metal1 s 14352 14790 14352 14790 4 _080_
rlabel metal1 s 16836 2550 16836 2550 4 _081_
rlabel metal1 s 15134 15674 15134 15674 4 _082_
rlabel metal1 s 15686 7820 15686 7820 4 _083_
rlabel metal2 s 1702 6205 1702 6205 4 _084_
rlabel metal2 s 16882 15980 16882 15980 4 _085_
rlabel metal3 s 6555 13260 6555 13260 4 _086_
rlabel metal1 s 15732 8058 15732 8058 4 _087_
rlabel metal2 s 18308 9588 18308 9588 4 _088_
rlabel metal2 s 15870 7990 15870 7990 4 _089_
rlabel metal1 s 18216 2618 18216 2618 4 _090_
rlabel metal1 s 9775 7922 9775 7922 4 _091_
rlabel metal1 s 3910 3570 3910 3570 4 _092_
rlabel metal3 s 17802 3179 17802 3179 4 _093_
rlabel metal1 s 5842 3162 5842 3162 4 _094_
rlabel metal2 s 12742 6766 12742 6766 4 _095_
rlabel metal1 s 14306 13294 14306 13294 4 _096_
rlabel metal1 s 2070 10778 2070 10778 4 _097_
rlabel metal1 s 11362 13294 11362 13294 4 _098_
rlabel metal1 s 8004 11798 8004 11798 4 _099_
rlabel metal1 s 13938 11118 13938 11118 4 _100_
rlabel metal1 s 4968 3502 4968 3502 4 _101_
rlabel metal1 s 3542 6664 3542 6664 4 _102_
rlabel metal1 s 15502 6086 15502 6086 4 _103_
rlabel metal1 s 2162 9962 2162 9962 4 _104_
rlabel metal1 s 2208 5882 2208 5882 4 _105_
rlabel metal2 s 16974 6477 16974 6477 4 _106_
rlabel metal3 s 5497 5508 5497 5508 4 _107_
rlabel metal1 s 1794 8364 1794 8364 4 _108_
rlabel metal1 s 14697 12818 14697 12818 4 _109_
rlabel metal1 s 6578 9146 6578 9146 4 _110_
rlabel metal1 s 5755 6358 5755 6358 4 _111_
rlabel metal1 s 4554 6222 4554 6222 4 _112_
rlabel metal1 s 5980 6154 5980 6154 4 _113_
rlabel metal2 s 8050 15011 8050 15011 4 _114_
rlabel metal2 s 14122 11016 14122 11016 4 _115_
rlabel metal1 s 12006 17204 12006 17204 4 _116_
rlabel metal3 s 13754 7259 13754 7259 4 _117_
rlabel metal1 s 16974 11594 16974 11594 4 _118_
rlabel metal1 s 18078 5338 18078 5338 4 _119_
rlabel metal3 s 14076 15504 14076 15504 4 _120_
rlabel metal2 s 1702 11900 1702 11900 4 _121_
rlabel metal1 s 14306 7922 14306 7922 4 _122_
rlabel metal2 s 15042 8109 15042 8109 4 _123_
rlabel metal1 s 1978 11730 1978 11730 4 _124_
rlabel metal2 s 3174 11832 3174 11832 4 _125_
rlabel metal1 s 6992 16626 6992 16626 4 _126_
rlabel metal1 s 5152 12070 5152 12070 4 _127_
rlabel metal1 s 18124 4590 18124 4590 4 _128_
rlabel metal1 s 17710 9588 17710 9588 4 _129_
rlabel metal4 s 17779 9588 17779 9588 4 _130_
rlabel metal2 s 18446 9078 18446 9078 4 _131_
rlabel metal2 s 12558 14620 12558 14620 4 _132_
rlabel metal2 s 12558 6171 12558 6171 4 _133_
rlabel metal1 s 10074 3026 10074 3026 4 _134_
rlabel metal1 s 10626 3060 10626 3060 4 _135_
rlabel metal3 s 10718 3043 10718 3043 4 _136_
rlabel metal2 s 10718 12274 10718 12274 4 _137_
rlabel metal1 s 12788 6358 12788 6358 4 _138_
rlabel metal2 s 17986 14195 17986 14195 4 _139_
rlabel metal1 s 13708 4794 13708 4794 4 _140_
rlabel metal1 s 16008 12886 16008 12886 4 _141_
rlabel metal1 s 7590 2482 7590 2482 4 _142_
rlabel metal2 s 15410 6171 15410 6171 4 _143_
rlabel metal3 s 16882 4675 16882 4675 4 _144_
rlabel metal2 s 2806 9180 2806 9180 4 _145_
rlabel metal1 s 7636 5678 7636 5678 4 _146_
rlabel metal2 s 4094 10455 4094 10455 4 _147_
rlabel metal2 s 15594 14433 15594 14433 4 _148_
rlabel metal3 s 14927 15436 14927 15436 4 _149_
rlabel metal1 s 9384 2618 9384 2618 4 _150_
rlabel metal3 s 4983 19788 4983 19788 4 clk
rlabel metal2 s 12834 10387 12834 10387 4 clknet_0_clk
rlabel metal1 s 1426 9418 1426 9418 4 clknet_2_0__leaf_clk
rlabel metal1 s 1978 12784 1978 12784 4 clknet_2_1__leaf_clk
rlabel metal1 s 12236 2482 12236 2482 4 clknet_2_2__leaf_clk
rlabel metal1 s 16422 9044 16422 9044 4 clknet_2_3__leaf_clk
rlabel metal2 s 12558 14076 12558 14076 4 net1
rlabel metal1 s 1610 13192 1610 13192 4 net10
rlabel metal1 s 2254 7752 2254 7752 4 net11
rlabel metal1 s 14214 14280 14214 14280 4 net12
rlabel metal2 s 1702 8381 1702 8381 4 net13
rlabel metal1 s 1564 2550 1564 2550 4 net14
rlabel metal1 s 1978 2618 1978 2618 4 net15
rlabel metal2 s 12558 4522 12558 4522 4 net16
rlabel metal1 s 6578 5610 6578 5610 4 net17
rlabel metal1 s 6095 2278 6095 2278 4 net18
rlabel metal1 s 14628 14926 14628 14926 4 net19
rlabel metal1 s 1610 8534 1610 8534 4 net2
rlabel metal1 s 14122 2822 14122 2822 4 net20
rlabel metal1 s 8050 2516 8050 2516 4 net21
rlabel metal1 s 11132 2618 11132 2618 4 net22
rlabel metal1 s 1886 16014 1886 16014 4 net23
rlabel metal1 s 1978 12206 1978 12206 4 net24
rlabel metal2 s 13846 13821 13846 13821 4 net25
rlabel metal1 s 3726 8534 3726 8534 4 net26
rlabel metal2 s 1886 7820 1886 7820 4 net27
rlabel metal2 s 1656 10132 1656 10132 4 net28
rlabel metal1 s 1886 5746 1886 5746 4 net29
rlabel metal1 s 1702 8466 1702 8466 4 net3
rlabel metal1 s 17986 9486 17986 9486 4 net30
rlabel metal3 s 13547 13804 13547 13804 4 net31
rlabel metal1 s 1886 3536 1886 3536 4 net32
rlabel metal1 s 1886 3060 1886 3060 4 net33
rlabel metal2 s 1886 2587 1886 2587 4 net34
rlabel metal1 s 12190 2992 12190 2992 4 net35
rlabel metal1 s 2668 9962 2668 9962 4 net36
rlabel metal1 s 5711 10710 5711 10710 4 net37
rlabel metal3 s 8648 8364 8648 8364 4 net38
rlabel metal2 s 13156 7684 13156 7684 4 net39
rlabel metal1 s 2944 8466 2944 8466 4 net4
rlabel metal2 s 11178 7616 11178 7616 4 net40
rlabel metal3 s 1326 9588 1326 9588 4 net41
rlabel metal3 s 1050 8908 1050 8908 4 net42
rlabel metal2 s 11822 11968 11822 11968 4 net5
rlabel metal1 s 17802 6800 17802 6800 4 net6
rlabel metal2 s 1610 14297 1610 14297 4 net7
rlabel metal2 s 1610 13991 1610 13991 4 net8
rlabel metal2 s 7130 10642 7130 10642 4 net9
rlabel metal1 s 1978 17204 1978 17204 4 rst_n
rlabel metal2 s 2714 17221 2714 17221 4 s_axi_araddr[0]
rlabel metal1 s 2898 17170 2898 17170 4 s_axi_araddr[1]
rlabel metal2 s 3082 17119 3082 17119 4 s_axi_araddr[2]
rlabel metal1 s 1472 17170 1472 17170 4 s_axi_araddr[3]
rlabel metal3 s 0 15648 800 15768 4 s_axi_arready
port 9 nsew
rlabel metal2 s 1426 15249 1426 15249 4 s_axi_arvalid
rlabel metal1 s 1334 14382 1334 14382 4 s_axi_awaddr[0]
rlabel metal2 s 1426 13787 1426 13787 4 s_axi_awaddr[1]
rlabel metal2 s 1978 13141 1978 13141 4 s_axi_awaddr[2]
rlabel metal1 s 1564 13294 1564 13294 4 s_axi_awaddr[3]
rlabel metal3 s 1142 11628 1142 11628 4 s_axi_awready
rlabel metal1 s 1748 11118 1748 11118 4 s_axi_awvalid
rlabel metal2 s 1426 10455 1426 10455 4 s_axi_bready
rlabel metal2 s 1610 8075 1610 8075 4 s_axi_bvalid
rlabel metal3 s 1418 7548 1418 7548 4 s_axi_rdata[0]
rlabel metal3 s 1142 6868 1142 6868 4 s_axi_rdata[1]
rlabel metal3 s 0 6128 800 6248 4 s_axi_rdata[2]
port 23 nsew
rlabel metal3 s 1142 5508 1142 5508 4 s_axi_rdata[3]
rlabel metal3 s 0 4768 800 4888 4 s_axi_rdata[4]
port 25 nsew
rlabel metal3 s 0 4088 800 4208 4 s_axi_rdata[5]
port 26 nsew
rlabel metal3 s 0 3408 800 3528 4 s_axi_rdata[6]
port 27 nsew
rlabel metal3 s 0 2728 800 2848 4 s_axi_rdata[7]
port 28 nsew
rlabel metal3 s 1418 2108 1418 2108 4 s_axi_rready
rlabel metal3 s 0 1368 800 1488 4 s_axi_rvalid
port 30 nsew
rlabel metal2 s 2806 1547 2806 1547 4 s_axi_wdata[0]
rlabel metal2 s 2898 1241 2898 1241 4 s_axi_wdata[1]
rlabel metal2 s 12282 1690 12282 1690 4 s_axi_wdata[2]
rlabel metal1 s 9752 2414 9752 2414 4 s_axi_wdata[3]
rlabel metal1 s 9108 2414 9108 2414 4 s_axi_wdata[4]
rlabel metal1 s 10396 2414 10396 2414 4 s_axi_wdata[5]
rlabel metal1 s 8648 2414 8648 2414 4 s_axi_wdata[6]
rlabel metal1 s 7728 2414 7728 2414 4 s_axi_wdata[7]
rlabel metal1 s 11776 2958 11776 2958 4 s_axi_wready
rlabel metal1 s 11178 2414 11178 2414 4 s_axi_wvalid
rlabel metal1 s 17618 11050 17618 11050 4 u_axi_slave.ctrl_reg\[0\]
rlabel metal1 s 7774 8602 7774 8602 4 u_axi_slave.ctrl_reg\[1\]
rlabel metal1 s 2208 12138 2208 12138 4 u_axi_slave.ctrl_reg\[2\]
rlabel metal1 s 6348 11322 6348 11322 4 u_axi_slave.ctrl_reg\[3\]
rlabel metal1 s 14444 9962 14444 9962 4 u_axi_slave.ctrl_reg\[4\]
rlabel metal3 s 3450 9571 3450 9571 4 u_axi_slave.ctrl_reg\[5\]
rlabel metal3 s 11362 11781 11362 11781 4 u_axi_slave.ctrl_reg\[6\]
rlabel metal2 s 14214 6035 14214 6035 4 u_axi_slave.ctrl_reg\[7\]
rlabel metal2 s 5704 6358 5704 6358 4 u_axi_slave.lfsr_data\[0\]
rlabel metal1 s 9522 16660 9522 16660 4 u_axi_slave.lfsr_data\[1\]
rlabel metal1 s 6900 7242 6900 7242 4 u_axi_slave.lfsr_data\[2\]
rlabel metal1 s 5336 7854 5336 7854 4 u_axi_slave.lfsr_data\[3\]
rlabel metal1 s 2254 6970 2254 6970 4 u_axi_slave.lfsr_data\[4\]
rlabel metal1 s 13478 2618 13478 2618 4 u_axi_slave.lfsr_data\[5\]
rlabel metal2 s 2162 6987 2162 6987 4 u_axi_slave.lfsr_data\[6\]
rlabel metal1 s 16376 13838 16376 13838 4 u_axi_slave.lfsr_data\[7\]
rlabel metal1 s 18768 2958 18768 2958 4 u_axi_slave.seed_reg\[0\]
rlabel metal2 s 9706 15198 9706 15198 4 u_axi_slave.seed_reg\[1\]
rlabel metal1 s 14168 8058 14168 8058 4 u_axi_slave.seed_reg\[2\]
rlabel metal1 s 6624 16082 6624 16082 4 u_axi_slave.seed_reg\[3\]
rlabel metal1 s 17940 8466 17940 8466 4 u_axi_slave.seed_reg\[4\]
rlabel metal1 s 14398 12920 14398 12920 4 u_axi_slave.seed_reg\[5\]
rlabel metal1 s 7590 6834 7590 6834 4 u_axi_slave.seed_reg\[6\]
rlabel metal1 s 6072 14586 6072 14586 4 u_axi_slave.seed_reg\[7\]
rlabel metal2 s 5060 13532 5060 13532 4 u_axi_slave.taps_reg\[0\]
rlabel metal2 s 6164 12988 6164 12988 4 u_axi_slave.taps_reg\[1\]
rlabel metal1 s 13616 11050 13616 11050 4 u_axi_slave.taps_reg\[2\]
rlabel metal1 s 18216 4114 18216 4114 4 u_axi_slave.taps_reg\[3\]
rlabel metal2 s 9614 8772 9614 8772 4 u_axi_slave.taps_reg\[4\]
rlabel metal1 s 9246 8908 9246 8908 4 u_axi_slave.taps_reg\[5\]
rlabel metal1 s 15180 15062 15180 15062 4 u_axi_slave.taps_reg\[6\]
rlabel metal1 s 7590 2278 7590 2278 4 u_axi_slave.taps_reg\[7\]
flabel metal5 s -1076 16004 21040 16324 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s -1076 12196 21040 12516 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s -1076 8388 21040 8708 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s -1076 4580 21040 4900 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 17140 -4 17460 19588 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 12701 -4 13021 19588 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8262 -4 8582 19588 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3823 -4 4143 19588 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 20720 -4 21040 19588 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s -1076 19268 21040 19588 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s -1076 -4 21040 316 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s -1076 -4 -756 19588 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s -1076 15344 21040 15664 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s -1076 11536 21040 11856 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s -1076 7728 21040 8048 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s -1076 3920 21040 4240 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 16480 -4 16800 19588 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12041 -4 12361 19588 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7602 -4 7922 19588 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3163 -4 3483 19588 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 20060 656 20380 18928 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal5 s -416 18608 20380 18928 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s -416 656 20380 976 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s -416 656 -96 18928 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 19728 800 19848 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 0 19048 800 19168 0 FreeSans 600 0 0 0 rst_n
port 4 nsew
flabel metal3 s 0 18368 800 18488 0 FreeSans 600 0 0 0 s_axi_araddr[0]
port 5 nsew
flabel metal3 s 0 17688 800 17808 0 FreeSans 600 0 0 0 s_axi_araddr[1]
port 6 nsew
flabel metal3 s 0 17008 800 17128 0 FreeSans 600 0 0 0 s_axi_araddr[2]
port 7 nsew
flabel metal3 s 0 16328 800 16448 0 FreeSans 600 0 0 0 s_axi_araddr[3]
port 8 nsew
flabel metal3 s 400 15708 400 15708 0 FreeSans 600 0 0 0 s_axi_arready
flabel metal3 s 0 14968 800 15088 0 FreeSans 600 0 0 0 s_axi_arvalid
port 10 nsew
flabel metal3 s 0 14288 800 14408 0 FreeSans 600 0 0 0 s_axi_awaddr[0]
port 11 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 s_axi_awaddr[1]
port 12 nsew
flabel metal3 s 0 12928 800 13048 0 FreeSans 600 0 0 0 s_axi_awaddr[2]
port 13 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 s_axi_awaddr[3]
port 14 nsew
flabel metal3 s 0 11568 800 11688 0 FreeSans 600 0 0 0 s_axi_awready
port 15 nsew
flabel metal3 s 0 10888 800 11008 0 FreeSans 600 0 0 0 s_axi_awvalid
port 16 nsew
flabel metal3 s 0 10208 800 10328 0 FreeSans 600 0 0 0 s_axi_bready
port 17 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 s_axi_bresp[0]
port 18 nsew
flabel metal3 s 0 8848 800 8968 0 FreeSans 600 0 0 0 s_axi_bresp[1]
port 19 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 s_axi_bvalid
port 20 nsew
flabel metal3 s 0 7488 800 7608 0 FreeSans 600 0 0 0 s_axi_rdata[0]
port 21 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 s_axi_rdata[1]
port 22 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 s_axi_rdata[2]
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 s_axi_rdata[3]
port 24 nsew
flabel metal3 s 400 4828 400 4828 0 FreeSans 600 0 0 0 s_axi_rdata[4]
flabel metal3 s 400 4148 400 4148 0 FreeSans 600 0 0 0 s_axi_rdata[5]
flabel metal3 s 400 3468 400 3468 0 FreeSans 600 0 0 0 s_axi_rdata[6]
flabel metal3 s 400 2788 400 2788 0 FreeSans 600 0 0 0 s_axi_rdata[7]
flabel metal3 s 0 2048 800 2168 0 FreeSans 600 0 0 0 s_axi_rready
port 29 nsew
flabel metal3 s 400 1428 400 1428 0 FreeSans 600 0 0 0 s_axi_rvalid
flabel metal3 s 0 688 800 808 0 FreeSans 600 0 0 0 s_axi_wdata[0]
port 31 nsew
flabel metal3 s 0 8 800 128 0 FreeSans 600 0 0 0 s_axi_wdata[1]
port 32 nsew
flabel metal2 s 12254 0 12310 800 0 FreeSans 280 90 0 0 s_axi_wdata[2]
port 33 nsew
flabel metal2 s 9678 0 9734 800 0 FreeSans 280 90 0 0 s_axi_wdata[3]
port 34 nsew
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 s_axi_wdata[4]
port 35 nsew
flabel metal2 s 10322 0 10378 800 0 FreeSans 280 90 0 0 s_axi_wdata[5]
port 36 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 s_axi_wdata[6]
port 37 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 s_axi_wdata[7]
port 38 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 s_axi_wready
port 39 nsew
flabel metal2 s 10966 0 11022 800 0 FreeSans 280 90 0 0 s_axi_wvalid
port 40 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
