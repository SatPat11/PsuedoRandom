* NGSPICE file created from lfsr_axi_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__lpflow_clkbufkapwr_1 abstract view
.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__lpflow_inputiso0n_1 abstract view
.subckt sky130_fd_sc_hd__lpflow_inputiso0n_1 A SLEEP_B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__lpflow_clkinvkapwr_1 abstract view
.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_1 A KAPWR VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_0 abstract view
.subckt sky130_fd_sc_hd__o21ai_0 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_0 abstract view
.subckt sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__lpflow_clkbufkapwr_4 abstract view
.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_4 A KAPWR VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__lpflow_isobufsrc_1 abstract view
.subckt sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__lpflow_clkbufkapwr_8 abstract view
.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_8 A KAPWR VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__lpflow_isobufsrc_4 abstract view
.subckt sky130_fd_sc_hd__lpflow_isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt lfsr_axi_top VGND VPWR clk rst_n s_axi_araddr[0] s_axi_araddr[1] s_axi_araddr[2]
+ s_axi_araddr[3] s_axi_arready s_axi_arvalid s_axi_awaddr[0] s_axi_awaddr[1] s_axi_awaddr[2]
+ s_axi_awaddr[3] s_axi_awready s_axi_awvalid s_axi_bready s_axi_bresp[0] s_axi_bresp[1]
+ s_axi_bvalid s_axi_rdata[0] s_axi_rdata[1] s_axi_rdata[2] s_axi_rdata[3] s_axi_rdata[4]
+ s_axi_rdata[5] s_axi_rdata[6] s_axi_rdata[7] s_axi_rready s_axi_rvalid s_axi_wdata[0]
+ s_axi_wdata[1] s_axi_wdata[2] s_axi_wdata[3] s_axi_wdata[4] s_axi_wdata[5] s_axi_wdata[6]
+ s_axi_wdata[7] s_axi_wready s_axi_wvalid
XANTENNA__203__B u_axi_slave.lfsr_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_294_ u_axi_slave.taps_reg\[4\] net18 _142_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__256__B1 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__340__RESET_B net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__247__B1 _112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_277_ _134_ _135_ _136_ _103_ net32 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__o32a_2
XANTENNA_fanout38_A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_200_ _071_ _072_ _073_ _074_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__o211a_2
XANTENNA__209__A u_axi_slave.lfsr_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_329_ clknet_2_0__leaf_clk _027_ net36 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__337__SET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input18_A s_axi_wdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__320__SET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__188__S _058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput31 net31 VGND VGND VPWR VPWR s_axi_rdata[5] sky130_fd_sc_hd__buf_4
XANTENNA__292__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__203__C u_axi_slave.taps_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_293_ _146_ _293_/KAPWR VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__265__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__256__B2 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__214__B _087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__247__A1 u_axi_slave.lfsr_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__247__B2 u_axi_slave.ctrl_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_276_ u_axi_slave.taps_reg\[6\] _107_ _112_ u_axi_slave.ctrl_reg\[6\] _114_ VGND
+ VGND VPWR VPWR _136_ sky130_fd_sc_hd__a221o_2
X_345_ clknet_2_1__leaf_clk _043_ net37 VGND VGND VPWR VPWR u_axi_slave.taps_reg\[7\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__257__SLEEP_B _112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__286__S _142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__174__A0 u_axi_slave.ctrl_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__209__B u_axi_slave.lfsr_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__156__A0 u_axi_slave.seed_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_328_ clknet_2_1__leaf_clk _026_ net37 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfrtp_2
XANTENNA__225__A u_axi_slave.lfsr_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_259_ _122_ _116_ _102_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output31_A net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__334__RESET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__294__S _142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__233__A u_axi_slave.lfsr_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput32 net32 VGND VGND VPWR VPWR s_axi_rdata[6] sky130_fd_sc_hd__buf_4
XANTENNA__283__A2 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__203__D u_axi_slave.taps_reg\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_292_ u_axi_slave.taps_reg\[3\] net17 _142_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__265__A2 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__247__A2 _111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_275_ u_axi_slave.lfsr_data\[6\] _111_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__lpflow_inputiso0n_1
XANTENNA__238__A2 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_344_ clknet_2_2__leaf_clk _042_ net38 VGND VGND VPWR VPWR u_axi_slave.taps_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__174__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__225__B _070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__241__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__209__C u_axi_slave.lfsr_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__156__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_327_ clknet_2_3__leaf_clk _025_ net40 VGND VGND VPWR VPWR u_axi_slave.lfsr_data\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_258_ u_axi_slave.taps_reg\[2\] _258_/KAPWR VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__lpflow_clkinvkapwr_1
X_189_ _066_ _189_/KAPWR VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__236__A _102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output24_A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__286__A0 u_axi_slave.taps_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__277__B1 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput33 net33 VGND VGND VPWR VPWR s_axi_rdata[7] sky130_fd_sc_hd__buf_4
XANTENNA__233__B _092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__259__B1 _102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_291_ _145_ _291_/KAPWR VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__244__A u_axi_slave.seed_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__256__A3 _120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__304__D _002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_343_ clknet_2_3__leaf_clk _041_ net39 VGND VGND VPWR VPWR u_axi_slave.taps_reg\[5\]
+ sky130_fd_sc_hd__dfstp_2
X_274_ u_axi_slave.seed_reg\[6\] _109_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__lpflow_inputiso0n_1
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__225__C _087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__209__D u_axi_slave.lfsr_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_188_ u_axi_slave.ctrl_reg\[7\] net21 _058_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__mux2_1
X_257_ u_axi_slave.ctrl_reg\[2\] _112_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__lpflow_inputiso0n_1
XANTENNA__151__B net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_326_ clknet_2_0__leaf_clk _024_ net36 VGND VGND VPWR VPWR u_axi_slave.lfsr_data\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_309_ clknet_2_1__leaf_clk _007_ net37 VGND VGND VPWR VPWR u_axi_slave.seed_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__286__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput23 net23 VGND VGND VPWR VPWR s_axi_arready sky130_fd_sc_hd__buf_4
Xoutput34 net34 VGND VGND VPWR VPWR s_axi_rvalid sky130_fd_sc_hd__buf_4
XANTENNA__277__B2 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input16_A s_axi_wdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A s_axi_awaddr[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_290_ u_axi_slave.taps_reg\[2\] net16 _142_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_342_ clknet_2_1__leaf_clk _040_ net38 VGND VGND VPWR VPWR u_axi_slave.taps_reg\[4\]
+ sky130_fd_sc_hd__dfstp_2
X_273_ net31 _103_ _132_ _133_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__o22a_2
XFILLER_0_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__235__SLEEP_B net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_256_ _117_ _119_ _120_ _103_ net27 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__o32a_2
XANTENNA__151__C net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ clknet_2_2__leaf_clk _023_ net39 VGND VGND VPWR VPWR u_axi_slave.lfsr_data\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_187_ _065_ _187_/KAPWR VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_308_ clknet_2_1__leaf_clk _006_ net37 VGND VGND VPWR VPWR u_axi_slave.seed_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_239_ _105_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__263__A u_axi_slave.lfsr_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__213__C1 _076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput24 net24 VGND VGND VPWR VPWR s_axi_awready sky130_fd_sc_hd__buf_4
XANTENNA__348__A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput35 net35 VGND VGND VPWR VPWR s_axi_wready sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__258__A u_axi_slave.taps_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__259__A2 _116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__318__D _016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__186__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_272_ u_axi_slave.seed_reg\[5\] _109_ _112_ u_axi_slave.ctrl_reg\[5\] _114_ VGND
+ VGND VPWR VPWR _133_ sky130_fd_sc_hd__a221o_2
XANTENNA__300__S _142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_341_ clknet_2_2__leaf_clk _039_ net40 VGND VGND VPWR VPWR u_axi_slave.taps_reg\[3\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__168__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__275__SLEEP_B _111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_255_ u_axi_slave.lfsr_data\[1\] _111_ _109_ u_axi_slave.seed_reg\[1\] VGND VGND
+ VPWR VPWR _120_ sky130_fd_sc_hd__a22o_2
X_186_ u_axi_slave.ctrl_reg\[6\] net20 _058_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_324_ clknet_2_2__leaf_clk _022_ net40 VGND VGND VPWR VPWR u_axi_slave.lfsr_data\[4\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload1 clknet_2_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_1
XPHY_EDGE_ROW_3_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_307_ clknet_2_3__leaf_clk _005_ net39 VGND VGND VPWR VPWR u_axi_slave.seed_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_169_ _055_ _169_/KAPWR VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XANTENNA__298__A0 u_axi_slave.taps_reg\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_238_ net34 _103_ _104_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__o21ai_0
XANTENNA__222__B1 _094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__204__B1 u_axi_slave.taps_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput25 net25 VGND VGND VPWR VPWR s_axi_bvalid sky130_fd_sc_hd__buf_4
XFILLER_0_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input21_A s_axi_wdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_271_ u_axi_slave.taps_reg\[5\] _107_ _111_ u_axi_slave.lfsr_data\[5\] VGND VGND
+ VPWR VPWR _132_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_340_ clknet_2_3__leaf_clk _038_ net1 VGND VGND VPWR VPWR u_axi_slave.taps_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__244__SLEEP_B _109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_323_ clknet_2_1__leaf_clk _021_ net37 VGND VGND VPWR VPWR u_axi_slave.lfsr_data\[3\]
+ sky130_fd_sc_hd__dfstp_4
X_185_ _064_ _185_/KAPWR VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XANTENNA__282__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_254_ _090_ _118_ _102_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o21ai_0
XANTENNA__192__A _068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload2 clknet_2_3__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_306_ clknet_2_1__leaf_clk _004_ net37 VGND VGND VPWR VPWR u_axi_slave.seed_reg\[4\]
+ sky130_fd_sc_hd__dfstp_2
X_237_ net13 net34 VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nand2_2
XANTENNA__298__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_168_ u_axi_slave.seed_reg\[6\] net20 _048_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__mux2_1
XANTENNA__222__B2 u_axi_slave.lfsr_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__222__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__213__A1 _081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__204__A1 u_axi_slave.lfsr_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__204__B2 u_axi_slave.lfsr_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput26 net26 VGND VGND VPWR VPWR s_axi_rdata[0] sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__198__B1 u_axi_slave.taps_reg\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A s_axi_wdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input6_A s_axi_arvalid VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__195__A u_axi_slave.ctrl_reg\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_270_ net30 _103_ _129_ _131_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__o22a_2
XFILLER_0_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ clknet_2_2__leaf_clk _020_ net39 VGND VGND VPWR VPWR u_axi_slave.lfsr_data\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_184_ u_axi_slave.ctrl_reg\[5\] net19 _058_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_253_ net5 _106_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__or2_0
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_305_ clknet_2_2__leaf_clk _003_ net39 VGND VGND VPWR VPWR u_axi_slave.seed_reg\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_167_ _054_ _167_/KAPWR VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
X_236_ _102_ _236_/KAPWR VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__lpflow_clkbufkapwr_4
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__213__A2 _082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_219_ u_axi_slave.lfsr_data\[0\] _070_ _089_ _093_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__204__A2 u_axi_slave.taps_reg\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput27 net27 VGND VGND VPWR VPWR s_axi_rdata[1] sky130_fd_sc_hd__buf_4
XANTENNA__198__B2 u_axi_slave.lfsr_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__198__A1 u_axi_slave.lfsr_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__195__B u_axi_slave.ctrl_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout40 net1 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_4
X_321_ clknet_2_0__leaf_clk _019_ net36 VGND VGND VPWR VPWR u_axi_slave.lfsr_data\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_183_ _063_ _183_/KAPWR VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__234__B1 _094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_252_ u_axi_slave.taps_reg\[1\] _116_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__lpflow_isobufsrc_1
XFILLER_0_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_235_ net23 net6 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__lpflow_inputiso0n_1
X_304_ clknet_2_0__leaf_clk _002_ net36 VGND VGND VPWR VPWR u_axi_slave.seed_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_166_ u_axi_slave.seed_reg\[5\] net19 _048_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_218_ _090_ u_axi_slave.seed_reg\[0\] _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__o21a_2
XFILLER_0_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput28 net28 VGND VGND VPWR VPWR s_axi_rdata[2] sky130_fd_sc_hd__buf_4
XFILLER_0_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__198__A2 u_axi_slave.taps_reg\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__264__D1 _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__270__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_182_ u_axi_slave.ctrl_reg\[4\] net18 _058_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__mux2_1
X_320_ clknet_2_3__leaf_clk _018_ net40 VGND VGND VPWR VPWR u_axi_slave.lfsr_data\[0\]
+ sky130_fd_sc_hd__dfstp_4
X_251_ net3 net2 net4 net5 VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__or4b_4
XFILLER_0_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__170__A0 u_axi_slave.seed_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__234__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__234__B2 u_axi_slave.lfsr_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__156__S _048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_165_ _053_ _165_/KAPWR VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XPHY_EDGE_ROW_23_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_303_ clknet_2_2__leaf_clk _001_ net39 VGND VGND VPWR VPWR u_axi_slave.seed_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_234_ _090_ u_axi_slave.seed_reg\[7\] _094_ u_axi_slave.lfsr_data\[6\] _101_ VGND
+ VGND VPWR VPWR _025_ sky130_fd_sc_hd__o221a_2
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_217_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__buf_4
Xoutput29 net29 VGND VGND VPWR VPWR s_axi_rdata[3] sky130_fd_sc_hd__buf_4
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__164__S _048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__270__A2 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__261__A2 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input12_A s_axi_bready VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input4_A s_axi_araddr[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_250_ net26 _103_ _115_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__o21ba_2
X_181_ _062_ _181_/KAPWR VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__170__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__234__A2 u_axi_slave.seed_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_302_ clknet_2_3__leaf_clk _000_ net40 VGND VGND VPWR VPWR u_axi_slave.seed_reg\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_233_ u_axi_slave.lfsr_data\[7\] _092_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__or2_0
XANTENNA__207__A2 _080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_164_ u_axi_slave.seed_reg\[4\] net18 _048_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__mux2_1
XANTENNA__279__SLEEP _116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_216_ u_axi_slave.ctrl_reg\[1\] u_axi_slave.ctrl_reg\[0\] VGND VGND VPWR VPWR _091_
+ sky130_fd_sc_hd__or2_0
XFILLER_0_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__180__S _058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__255__B1 _109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__228__B1 _092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_180_ u_axi_slave.ctrl_reg\[3\] net17 _058_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__219__B1 _089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_232_ _090_ u_axi_slave.seed_reg\[6\] _094_ u_axi_slave.lfsr_data\[5\] _100_ VGND
+ VGND VPWR VPWR _024_ sky130_fd_sc_hd__o221a_2
X_163_ _052_ _163_/KAPWR VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_301_ _150_ _301_/KAPWR VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_215_ _086_ _215_/KAPWR VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__lpflow_clkbufkapwr_8
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__178__S _058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__273__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__255__A1 u_axi_slave.lfsr_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__249__D1 _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__220__A _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__228__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__228__B2 u_axi_slave.lfsr_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__186__S _058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__219__B2 _093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__219__A1 u_axi_slave.lfsr_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__164__A0 u_axi_slave.seed_reg\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_162_ u_axi_slave.seed_reg\[3\] net17 _048_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__mux2_1
X_231_ u_axi_slave.lfsr_data\[6\] _092_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__or2_0
X_300_ u_axi_slave.taps_reg\[7\] net21 _142_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__300__A0 u_axi_slave.taps_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output29_A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput1 rst_n VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_214_ _083_ _087_ _088_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__223__A u_axi_slave.lfsr_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__276__C1 _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__273__A2 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__264__A2 _112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__255__A2 _111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__191__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__182__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__220__B u_axi_slave.ctrl_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__228__A2 u_axi_slave.seed_reg\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__292__S _142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__219__A2 _070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input10_A s_axi_awaddr[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__231__A u_axi_slave.lfsr_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__164__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__268__SLEEP _116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input2_A s_axi_araddr[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_161_ _051_ _161_/KAPWR VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_230_ _090_ u_axi_slave.seed_reg\[5\] _094_ u_axi_slave.lfsr_data\[4\] _099_ VGND
+ VGND VPWR VPWR _023_ sky130_fd_sc_hd__o221a_2
XFILLER_0_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 s_axi_araddr[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__300__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_213_ _081_ _082_ _075_ _076_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__a211o_2
XFILLER_0_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__294__A0 u_axi_slave.taps_reg\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__223__B _092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__276__B1 _112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__267__B1 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__191__A2 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__327__RESET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__229__A u_axi_slave.lfsr_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__231__B _092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_160_ u_axi_slave.seed_reg\[2\] net16 _048_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 s_axi_araddr[1] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__298__S _142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_289_ _144_ _289_/KAPWR VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
X_212_ _084_ _085_ _086_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__294__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__276__A1 u_axi_slave.taps_reg\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__249__A1 u_axi_slave.taps_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__176__A0 u_axi_slave.ctrl_reg\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__229__B _092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__245__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout36 net38 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_4
XFILLER_0_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 s_axi_araddr[2] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_288_ u_axi_slave.taps_reg\[1\] net15 _142_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_211_ u_axi_slave.ctrl_reg\[1\] _211_/KAPWR VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__lpflow_clkinvkapwr_1
XFILLER_0_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output27_A net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__253__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__276__A2 _107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__248__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__194__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__249__A2 _107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__274__SLEEP_B _109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__176__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__158__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout37 net38 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_18_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__171__A _056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__316__D _014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 s_axi_araddr[3] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_0_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__230__B1 _094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_287_ _143_ _287_/KAPWR VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
X_210_ u_axi_slave.lfsr_data\[1\] u_axi_slave.lfsr_data\[0\] u_axi_slave.lfsr_data\[3\]
+ u_axi_slave.lfsr_data\[2\] VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__or4_2
XFILLER_0_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout39_A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__253__B _106_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_339_ clknet_2_3__leaf_clk _037_ net1 VGND VGND VPWR VPWR u_axi_slave.taps_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__248__B net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__194__A2 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input19_A s_axi_wdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__319__D _017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout38 net1 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_4_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__230__B2 u_axi_slave.lfsr_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__230__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_286_ u_axi_slave.taps_reg\[0\] net14 _142_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__mux2_1
Xinput6 s_axi_arvalid VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XANTENNA__327__D _025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__288__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ clknet_2_1__leaf_clk _036_ net37 VGND VGND VPWR VPWR u_axi_slave.taps_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ u_axi_slave.lfsr_data\[4\] _111_ _109_ u_axi_slave.seed_reg\[4\] _130_ VGND
+ VGND VPWR VPWR _131_ sky130_fd_sc_hd__a221o_2
XFILLER_0_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput20 s_axi_wdata[6] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XANTENNA_output32_A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__340__D _038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__190__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__275__A u_axi_slave.lfsr_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__335__D _033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout39 net40 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_4
XFILLER_0_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_285_ _141_ _285_/KAPWR VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__lpflow_clkbufkapwr_4
Xinput7 s_axi_awaddr[0] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XANTENNA__206__C1 _080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_268_ u_axi_slave.taps_reg\[4\] _116_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__lpflow_isobufsrc_1
X_199_ u_axi_slave.lfsr_data\[5\] u_axi_slave.lfsr_data\[4\] u_axi_slave.taps_reg\[4\]
+ u_axi_slave.taps_reg\[5\] VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__nand4_4
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_337_ clknet_2_2__leaf_clk _035_ net40 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfstp_4
XTAP_TAPCELL_ROW_11_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__188__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__197__A1 u_axi_slave.lfsr_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__197__B2 u_axi_slave.lfsr_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output25_A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 s_axi_awaddr[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
Xinput21 s_axi_wdata[7] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__260__B1 _109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__314__RESET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__196__A u_axi_slave.lfsr_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__224__B1 _094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_284_ net9 net10 _044_ _046_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__and4b_2
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput8 s_axi_awaddr[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_336_ clknet_2_3__leaf_clk _034_ net38 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfrtp_2
X_267_ _128_ _118_ _103_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__o21ai_0
X_198_ u_axi_slave.lfsr_data\[4\] u_axi_slave.taps_reg\[4\] u_axi_slave.taps_reg\[5\]
+ u_axi_slave.lfsr_data\[5\] VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__339__RESET_B net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__197__A2 u_axi_slave.taps_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__289__A _144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput11 s_axi_awvalid VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XANTENNA__199__A u_axi_slave.lfsr_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput22 s_axi_wvalid VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
X_319_ clknet_2_0__leaf_clk _017_ net36 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfstp_2
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__193__B1_N net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__252__SLEEP _116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__260__A1 u_axi_slave.lfsr_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__260__B2 u_axi_slave.seed_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input17_A s_axi_wdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__196__B u_axi_slave.lfsr_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input9_A s_axi_awaddr[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__224__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__224__B2 u_axi_slave.lfsr_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__160__A0 u_axi_slave.seed_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 s_axi_awaddr[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_0_11_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_283_ _140_ net6 _104_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_1_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_335_ clknet_2_1__leaf_clk _033_ net37 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfrtp_2
X_197_ u_axi_slave.lfsr_data\[0\] u_axi_slave.taps_reg\[0\] u_axi_slave.taps_reg\[1\]
+ u_axi_slave.lfsr_data\[1\] VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__a22oi_4
X_266_ u_axi_slave.ctrl_reg\[4\] _266_/KAPWR VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__lpflow_clkinvkapwr_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput12 s_axi_bready VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
X_249_ u_axi_slave.taps_reg\[0\] _107_ _110_ _113_ _114_ VGND VGND VPWR VPWR _115_
+ sky130_fd_sc_hd__a2111oi_2
XANTENNA__199__B u_axi_slave.lfsr_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_318_ clknet_2_0__leaf_clk _016_ net36 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__272__C1 _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output30_A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__260__A2 _111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__196__C u_axi_slave.taps_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__162__S _048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__224__A2 u_axi_slave.seed_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__160__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_282_ net23 VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__inv_2
X_334_ clknet_2_3__leaf_clk _032_ net40 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_265_ net29 _103_ _127_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__o21ba_2
X_196_ u_axi_slave.lfsr_data\[1\] u_axi_slave.lfsr_data\[0\] u_axi_slave.taps_reg\[0\]
+ u_axi_slave.taps_reg\[1\] VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__and4_2
XFILLER_0_2_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__290__A0 u_axi_slave.taps_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_179_ _061_ _179_/KAPWR VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
X_248_ net23 net6 VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__nand2_4
Xinput13 s_axi_rready VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_317_ clknet_2_2__leaf_clk _015_ net39 VGND VGND VPWR VPWR u_axi_slave.ctrl_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__170__S _048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__199__C u_axi_slave.taps_reg\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__272__B1 _112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_output23_A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__254__B1 _102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A s_axi_wvalid VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__218__B1 _092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_281_ net33 _103_ _139_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_264_ u_axi_slave.ctrl_reg\[3\] _112_ _125_ _126_ _114_ VGND VGND VPWR VPWR _127_
+ sky130_fd_sc_hd__a2111oi_2
X_195_ u_axi_slave.ctrl_reg\[1\] u_axi_slave.ctrl_reg\[0\] VGND VGND VPWR VPWR _070_
+ sky130_fd_sc_hd__nor2_2
XFILLER_0_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ clknet_2_2__leaf_clk _031_ net36 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfrtp_2
XANTENNA__241__SLEEP _106_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__168__S _048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_316_ clknet_2_3__leaf_clk _014_ net40 VGND VGND VPWR VPWR u_axi_slave.ctrl_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__290__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput14 s_axi_wdata[0] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
X_247_ u_axi_slave.lfsr_data\[0\] _111_ _112_ u_axi_slave.ctrl_reg\[0\] VGND VGND
+ VPWR VPWR _113_ sky130_fd_sc_hd__a22o_2
XANTENNA__281__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__199__D u_axi_slave.taps_reg\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_178_ u_axi_slave.ctrl_reg\[2\] net16 _058_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__mux2_1
XANTENNA__272__B2 u_axi_slave.ctrl_reg\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__210__A u_axi_slave.lfsr_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__254__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__176__S _058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__205__A u_axi_slave.lfsr_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input15_A s_axi_wdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__218__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_280_ u_axi_slave.ctrl_reg\[7\] _112_ _137_ _138_ _114_ VGND VGND VPWR VPWR _139_
+ sky130_fd_sc_hd__a2111oi_2
XANTENNA_input7_A s_axi_awaddr[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_263_ u_axi_slave.lfsr_data\[3\] _111_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__lpflow_inputiso0n_1
X_194_ net12 net25 _069_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a21o_2
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_332_ clknet_2_2__leaf_clk _030_ net36 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__184__S _058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_246_ net5 _106_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__nor2_4
X_177_ _060_ _177_/KAPWR VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XANTENNA__281__A2 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_315_ clknet_2_0__leaf_clk _013_ net36 VGND VGND VPWR VPWR u_axi_slave.ctrl_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput15 s_axi_wdata[1] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XANTENNA__272__A2 _109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_229_ u_axi_slave.lfsr_data\[5\] _092_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__or2_0
XFILLER_0_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__210__B u_axi_slave.lfsr_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__205__B u_axi_slave.lfsr_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__221__A u_axi_slave.lfsr_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__218__A2 u_axi_slave.seed_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__216__A u_axi_slave.ctrl_reg\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_262_ u_axi_slave.taps_reg\[3\] _107_ _109_ u_axi_slave.seed_reg\[3\] VGND VGND VPWR
+ VPWR _125_ sky130_fd_sc_hd__a22o_2
X_331_ clknet_2_0__leaf_clk _029_ net36 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_4
X_193_ net22 net11 net24 VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__a21boi_2
XANTENNA__290__S _142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__341__SET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_176_ u_axi_slave.ctrl_reg\[1\] net15 _058_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__mux2_1
X_245_ net5 _108_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__lpflow_isobufsrc_4
X_314_ clknet_2_3__leaf_clk _012_ net40 VGND VGND VPWR VPWR u_axi_slave.ctrl_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput16 s_axi_wdata[2] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_228_ _090_ u_axi_slave.seed_reg\[4\] _092_ u_axi_slave.lfsr_data\[4\] _098_ VGND
+ VGND VPWR VPWR _022_ sky130_fd_sc_hd__o221a_2
X_159_ _050_ _159_/KAPWR VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XANTENNA__210__C u_axi_slave.lfsr_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout40_A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__205__C u_axi_slave.taps_reg\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__221__B _092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__216__B u_axi_slave.ctrl_reg\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input20_A s_axi_wdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__288__S _142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_192_ _068_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__buf_1
XANTENNA__227__A u_axi_slave.lfsr_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_261_ net28 _103_ _121_ _124_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__o22a_2
XFILLER_0_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_330_ clknet_2_2__leaf_clk _028_ net39 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_313_ clknet_2_1__leaf_clk _011_ net37 VGND VGND VPWR VPWR u_axi_slave.ctrl_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_16_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_175_ _059_ _175_/KAPWR VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
X_244_ u_axi_slave.seed_reg\[0\] _109_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__lpflow_inputiso0n_1
Xinput17 s_axi_wdata[3] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__184__A0 u_axi_slave.ctrl_reg\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_227_ u_axi_slave.lfsr_data\[3\] _070_ _087_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__or3_2
XANTENNA__296__S _142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_158_ u_axi_slave.seed_reg\[1\] net15 _048_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__mux2_1
XANTENNA__210__D u_axi_slave.lfsr_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__235__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__205__D u_axi_slave.taps_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__324__SET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input13_A s_axi_rready VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ u_axi_slave.lfsr_data\[2\] _111_ _109_ u_axi_slave.seed_reg\[2\] _123_ VGND
+ VGND VPWR VPWR _124_ sky130_fd_sc_hd__a221o_2
XANTENNA_input5_A s_axi_araddr[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__227__B _070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__243__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_191_ net12 net25 _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__a21boi_2
X_174_ u_axi_slave.ctrl_reg\[0\] net14 _058_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__mux2_1
X_243_ net5 _108_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_16_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 s_axi_wdata[4] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
X_312_ clknet_2_2__leaf_clk _010_ net39 VGND VGND VPWR VPWR u_axi_slave.ctrl_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_21_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__184__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_226_ _090_ u_axi_slave.seed_reg\[3\] _092_ u_axi_slave.lfsr_data\[3\] _097_ VGND
+ VGND VPWR VPWR _021_ sky130_fd_sc_hd__o221a_2
X_157_ _049_ _157_/KAPWR VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XANTENNA__166__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_209_ u_axi_slave.lfsr_data\[5\] u_axi_slave.lfsr_data\[4\] u_axi_slave.lfsr_data\[7\]
+ u_axi_slave.lfsr_data\[6\] VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__or4_2
XANTENNA__246__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__296__A0 u_axi_slave.taps_reg\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__227__C _087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__278__B1 _109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_190_ net25 _044_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__or2_0
XANTENNA__202__B1 u_axi_slave.taps_reg\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__269__B1 _109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_173_ _057_ _173_/KAPWR VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__lpflow_clkbufkapwr_4
X_311_ clknet_2_1__leaf_clk _009_ net37 VGND VGND VPWR VPWR u_axi_slave.ctrl_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_16_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ net3 net2 net4 VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__or3b_4
Xinput19 s_axi_wdata[5] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__193__A2 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_156_ u_axi_slave.seed_reg\[0\] net14 _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__mux2_1
X_225_ u_axi_slave.lfsr_data\[2\] _070_ _087_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_9_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_208_ _075_ _076_ _081_ _082_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__o211a_2
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__246__B _106_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__257__A u_axi_slave.ctrl_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__296__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__278__B2 u_axi_slave.seed_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__278__A1 u_axi_slave.lfsr_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__202__A1 u_axi_slave.lfsr_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__202__B2 u_axi_slave.lfsr_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__269__B2 u_axi_slave.seed_reg\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__269__A1 u_axi_slave.lfsr_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ clknet_2_3__leaf_clk _008_ net39 VGND VGND VPWR VPWR u_axi_slave.ctrl_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_172_ net9 _045_ _046_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__and3b_2
X_241_ net5 _106_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__lpflow_isobufsrc_4
XTAP_TAPCELL_ROW_21_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__178__A0 u_axi_slave.ctrl_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_224_ _090_ u_axi_slave.seed_reg\[2\] _094_ u_axi_slave.lfsr_data\[1\] _096_ VGND
+ VGND VPWR VPWR _020_ sky130_fd_sc_hd__o221a_2
X_155_ _047_ _155_/KAPWR VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__lpflow_clkbufkapwr_4
XPHY_EDGE_ROW_25_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_207_ _079_ _080_ _077_ _078_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__278__A2 _111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__268__A u_axi_slave.taps_reg\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__202__A2 u_axi_slave.taps_reg\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input11_A s_axi_awvalid VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__269__A2 _111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input3_A s_axi_araddr[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_240_ net3 net2 net4 VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__or3_4
X_171_ _056_ _171_/KAPWR VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__178__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_223_ u_axi_slave.lfsr_data\[2\] _092_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__or2_0
XFILLER_0_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_154_ net9 _045_ _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__and3_2
Xlfsr_axi_top_41 VGND VGND VPWR VPWR lfsr_axi_top_41/HI s_axi_bresp[0] sky130_fd_sc_hd__conb_1
XFILLER_0_20_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_206_ _077_ _078_ _079_ _080_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__a211o_2
XFILLER_0_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__232__B1 _094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__251__D_N net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__152__SLEEP net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_170_ u_axi_slave.seed_reg\[7\] net21 _048_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__mux2_2
XANTENNA__279__A u_axi_slave.taps_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_299_ _149_ _299_/KAPWR VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__280__D1 _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_222_ _090_ u_axi_slave.seed_reg\[1\] _094_ u_axi_slave.lfsr_data\[0\] _095_ VGND
+ VGND VPWR VPWR _019_ sky130_fd_sc_hd__o221a_2
X_153_ net8 net7 VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__nor2_2
Xlfsr_axi_top_42 VGND VGND VPWR VPWR lfsr_axi_top_42/HI s_axi_bresp[1] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_8_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_205_ u_axi_slave.lfsr_data\[7\] u_axi_slave.lfsr_data\[6\] u_axi_slave.taps_reg\[6\]
+ u_axi_slave.taps_reg\[7\] VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__and4_2
XFILLER_0_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__232__B2 u_axi_slave.lfsr_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__232__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__284__B net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_298_ u_axi_slave.taps_reg\[6\] net20 _142_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__mux2_1
XANTENNA__302__SET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_221_ u_axi_slave.lfsr_data\[1\] _092_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__or2_0
X_152_ _044_ net10 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__lpflow_isobufsrc_1
XTAP_TAPCELL_ROW_8_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_204_ u_axi_slave.lfsr_data\[6\] u_axi_slave.taps_reg\[6\] u_axi_slave.taps_reg\[7\]
+ u_axi_slave.lfsr_data\[7\] VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a22oi_4
XANTENNA__250__A2 _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__208__C1 _082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 _024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_297_ _148_ _297_/KAPWR VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XFILLER_0_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__160__S _048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__271__B1 _111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input1_A rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_151_ net22 net11 net24 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__and3_2
X_220_ _090_ u_axi_slave.ctrl_reg\[0\] VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__nand2_4
XANTENNA__262__B1 _109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_203_ u_axi_slave.lfsr_data\[3\] u_axi_slave.lfsr_data\[2\] u_axi_slave.taps_reg\[2\]
+ u_axi_slave.taps_reg\[3\] VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__nand4_4
XPHY_EDGE_ROW_4_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__226__B1 _092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__208__B1 _081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__316__RESET_B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__158__S _048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_296_ u_axi_slave.taps_reg\[5\] net19 _142_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__271__B2 u_axi_slave.lfsr_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__271__A1 u_axi_slave.taps_reg\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__262__A1 u_axi_slave.taps_reg\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ net24 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
X_279_ u_axi_slave.taps_reg\[7\] _116_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__lpflow_isobufsrc_1
X_202_ u_axi_slave.lfsr_data\[2\] u_axi_slave.taps_reg\[2\] u_axi_slave.taps_reg\[3\]
+ u_axi_slave.lfsr_data\[3\] VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__a22o_2
XANTENNA__226__A1 _090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__226__B2 u_axi_slave.lfsr_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output33_A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__166__S _048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__174__S _058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__203__A u_axi_slave.lfsr_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_295_ _147_ _295_/KAPWR VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__lpflow_clkbufkapwr_1
XANTENNA__280__A2 _112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__271__A2 _107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__262__A2 _107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_278_ u_axi_slave.lfsr_data\[7\] _111_ _109_ u_axi_slave.seed_reg\[7\] VGND VGND
+ VPWR VPWR _137_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__180__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_201_ _073_ _074_ _071_ _072_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_19_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__162__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__182__S _058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__211__A u_axi_slave.ctrl_reg\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__208__A2 _076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__263__SLEEP_B _111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput30 net30 VGND VGND VPWR VPWR s_axi_rdata[4] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_18_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__292__A0 u_axi_slave.taps_reg\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

